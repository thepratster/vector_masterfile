-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity vector_control_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity vector_control_daemon;
architecture Default of vector_control_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal vector_control_daemon_CP_8401_start: Boolean;
  signal vector_control_daemon_CP_8401_symbol: Boolean;
  -- links between control-path and data-path
  signal MUL_f32_f32_1916_inst_ack_0 : boolean;
  signal if_stmt_1962_branch_ack_1 : boolean;
  signal if_stmt_1962_branch_ack_0 : boolean;
  signal if_stmt_1962_branch_req_0 : boolean;
  signal EQ_f32_u1_1960_inst_req_0 : boolean;
  signal EQ_f32_u1_1960_inst_req_1 : boolean;
  signal ADD_f32_f32_1940_inst_req_0 : boolean;
  signal SHL_u32_u32_1997_inst_req_0 : boolean;
  signal SHL_u32_u32_1997_inst_ack_0 : boolean;
  signal EQ_f32_u1_1960_inst_ack_0 : boolean;
  signal AND_u32_u32_1979_inst_req_1 : boolean;
  signal AND_u32_u32_1979_inst_ack_1 : boolean;
  signal AND_u32_u32_1979_inst_req_0 : boolean;
  signal AND_u32_u32_1979_inst_ack_0 : boolean;
  signal EQ_f32_u1_1960_inst_ack_1 : boolean;
  signal XOR_u32_u32_2312_inst_ack_1 : boolean;
  signal SHL_u32_u32_1997_inst_req_1 : boolean;
  signal SHL_u32_u32_1997_inst_ack_1 : boolean;
  signal SUB_u32_u32_2322_inst_ack_0 : boolean;
  signal LSHR_u32_u32_1985_inst_req_1 : boolean;
  signal LSHR_u32_u32_1985_inst_ack_1 : boolean;
  signal AND_u32_u32_1991_inst_req_0 : boolean;
  signal AND_u32_u32_1991_inst_ack_0 : boolean;
  signal type_cast_1954_inst_req_0 : boolean;
  signal type_cast_1954_inst_ack_0 : boolean;
  signal AND_u32_u32_1991_inst_req_1 : boolean;
  signal AND_u32_u32_1991_inst_ack_1 : boolean;
  signal MUL_f32_f32_1916_inst_req_0 : boolean;
  signal LSHR_u32_u32_1985_inst_req_0 : boolean;
  signal LSHR_u32_u32_1985_inst_ack_0 : boolean;
  signal RPIPE_in_data_1720_inst_req_0 : boolean;
  signal RPIPE_in_data_1720_inst_ack_0 : boolean;
  signal RPIPE_in_data_1720_inst_req_1 : boolean;
  signal RPIPE_in_data_1720_inst_ack_1 : boolean;
  signal RPIPE_in_data_1723_inst_req_0 : boolean;
  signal RPIPE_in_data_1723_inst_ack_0 : boolean;
  signal RPIPE_in_data_1723_inst_req_1 : boolean;
  signal RPIPE_in_data_1723_inst_ack_1 : boolean;
  signal RPIPE_in_data_1726_inst_req_0 : boolean;
  signal RPIPE_in_data_1726_inst_ack_0 : boolean;
  signal RPIPE_in_data_1726_inst_req_1 : boolean;
  signal RPIPE_in_data_1726_inst_ack_1 : boolean;
  signal RPIPE_in_data_1729_inst_req_0 : boolean;
  signal RPIPE_in_data_1729_inst_ack_0 : boolean;
  signal RPIPE_in_data_1729_inst_req_1 : boolean;
  signal RPIPE_in_data_1729_inst_ack_1 : boolean;
  signal RPIPE_in_data_1732_inst_req_0 : boolean;
  signal RPIPE_in_data_1732_inst_ack_0 : boolean;
  signal RPIPE_in_data_1732_inst_req_1 : boolean;
  signal RPIPE_in_data_1732_inst_ack_1 : boolean;
  signal SLT_f32_u1_1737_inst_req_0 : boolean;
  signal SLT_f32_u1_1737_inst_ack_0 : boolean;
  signal SLT_f32_u1_1737_inst_req_1 : boolean;
  signal SLT_f32_u1_1737_inst_ack_1 : boolean;
  signal if_stmt_1739_branch_req_0 : boolean;
  signal if_stmt_1739_branch_ack_1 : boolean;
  signal if_stmt_1739_branch_ack_0 : boolean;
  signal type_cast_1749_inst_req_0 : boolean;
  signal type_cast_1749_inst_ack_0 : boolean;
  signal type_cast_1749_inst_req_1 : boolean;
  signal type_cast_1749_inst_ack_1 : boolean;
  signal ADD_f64_f64_1755_inst_req_0 : boolean;
  signal ADD_f64_f64_1755_inst_ack_0 : boolean;
  signal ADD_f64_f64_1755_inst_req_1 : boolean;
  signal ADD_f64_f64_1755_inst_ack_1 : boolean;
  signal type_cast_1759_inst_req_0 : boolean;
  signal type_cast_1759_inst_ack_0 : boolean;
  signal type_cast_1759_inst_req_1 : boolean;
  signal type_cast_1759_inst_ack_1 : boolean;
  signal SGT_f32_u1_1766_inst_req_0 : boolean;
  signal SGT_f32_u1_1766_inst_ack_0 : boolean;
  signal SGT_f32_u1_1766_inst_req_1 : boolean;
  signal SGT_f32_u1_1766_inst_ack_1 : boolean;
  signal if_stmt_1768_branch_req_0 : boolean;
  signal if_stmt_1768_branch_ack_1 : boolean;
  signal if_stmt_1768_branch_ack_0 : boolean;
  signal type_cast_1777_inst_req_0 : boolean;
  signal type_cast_1777_inst_ack_0 : boolean;
  signal type_cast_1777_inst_req_1 : boolean;
  signal type_cast_1777_inst_ack_1 : boolean;
  signal ADD_f64_f64_1783_inst_req_0 : boolean;
  signal ADD_f64_f64_1783_inst_ack_0 : boolean;
  signal ADD_f64_f64_1783_inst_req_1 : boolean;
  signal ADD_f64_f64_1783_inst_ack_1 : boolean;
  signal type_cast_1787_inst_req_0 : boolean;
  signal type_cast_1787_inst_ack_0 : boolean;
  signal type_cast_1787_inst_req_1 : boolean;
  signal type_cast_1787_inst_ack_1 : boolean;
  signal if_stmt_1905_branch_req_0 : boolean;
  signal MUL_f32_f32_1804_inst_req_0 : boolean;
  signal MUL_f32_f32_1804_inst_ack_0 : boolean;
  signal MUL_f32_f32_1804_inst_req_1 : boolean;
  signal MUL_f32_f32_1804_inst_ack_1 : boolean;
  signal MUL_f32_f32_1916_inst_ack_1 : boolean;
  signal LSHR_u32_u32_1973_inst_ack_1 : boolean;
  signal SGT_f32_u1_1903_inst_ack_1 : boolean;
  signal MUL_f32_f32_1935_inst_ack_1 : boolean;
  signal MUL_f32_f32_1916_inst_req_1 : boolean;
  signal type_cast_1950_inst_ack_1 : boolean;
  signal MUL_f32_f32_1935_inst_req_1 : boolean;
  signal SGT_f32_u1_1903_inst_req_1 : boolean;
  signal ADD_f32_f32_1809_inst_req_0 : boolean;
  signal ADD_f32_f32_1809_inst_ack_0 : boolean;
  signal ADD_f32_f32_1809_inst_req_1 : boolean;
  signal ADD_f32_f32_1809_inst_ack_1 : boolean;
  signal LSHR_u32_u32_1973_inst_req_1 : boolean;
  signal XOR_u32_u32_2312_inst_req_1 : boolean;
  signal type_cast_1950_inst_req_1 : boolean;
  signal if_stmt_1905_branch_ack_0 : boolean;
  signal SGT_f32_u1_1903_inst_ack_0 : boolean;
  signal MUL_f32_f32_1946_inst_ack_1 : boolean;
  signal MUL_f32_f32_1946_inst_req_1 : boolean;
  signal SGT_f32_u1_1903_inst_req_0 : boolean;
  signal SUB_f32_f32_1814_inst_req_0 : boolean;
  signal SUB_f32_f32_1814_inst_ack_0 : boolean;
  signal SUB_f32_f32_1814_inst_req_1 : boolean;
  signal SUB_f32_f32_1814_inst_ack_1 : boolean;
  signal MUL_f32_f32_1946_inst_ack_0 : boolean;
  signal MUL_f32_f32_1946_inst_req_0 : boolean;
  signal type_cast_1950_inst_ack_0 : boolean;
  signal ADD_f32_f32_1819_inst_req_0 : boolean;
  signal ADD_f32_f32_1819_inst_ack_0 : boolean;
  signal ADD_f32_f32_1819_inst_req_1 : boolean;
  signal ADD_f32_f32_1819_inst_ack_1 : boolean;
  signal LSHR_u32_u32_1973_inst_req_0 : boolean;
  signal LSHR_u32_u32_1973_inst_ack_0 : boolean;
  signal MUL_f32_f32_1935_inst_ack_0 : boolean;
  signal MUL_f32_f32_1825_inst_req_0 : boolean;
  signal MUL_f32_f32_1825_inst_ack_0 : boolean;
  signal MUL_f32_f32_1825_inst_req_1 : boolean;
  signal MUL_f32_f32_1825_inst_ack_1 : boolean;
  signal if_stmt_1892_branch_ack_0 : boolean;
  signal MUL_f32_f32_1935_inst_req_0 : boolean;
  signal type_cast_1950_inst_req_0 : boolean;
  signal ADD_f32_f32_1830_inst_req_0 : boolean;
  signal ADD_f32_f32_1830_inst_ack_0 : boolean;
  signal ADD_f32_f32_1830_inst_req_1 : boolean;
  signal ADD_f32_f32_1830_inst_ack_1 : boolean;
  signal ADD_f32_f32_1940_inst_ack_1 : boolean;
  signal ADD_f32_f32_1940_inst_req_1 : boolean;
  signal if_stmt_1892_branch_ack_1 : boolean;
  signal if_stmt_1892_branch_req_0 : boolean;
  signal type_cast_1834_inst_req_0 : boolean;
  signal type_cast_1834_inst_ack_0 : boolean;
  signal type_cast_1834_inst_req_1 : boolean;
  signal type_cast_1834_inst_ack_1 : boolean;
  signal ADD_f32_f32_1940_inst_ack_0 : boolean;
  signal if_stmt_1905_branch_ack_1 : boolean;
  signal SLT_f64_u1_1840_inst_req_0 : boolean;
  signal SLT_f64_u1_1840_inst_ack_0 : boolean;
  signal SLT_f32_u1_1890_inst_ack_1 : boolean;
  signal SLT_f64_u1_1840_inst_req_1 : boolean;
  signal SLT_f64_u1_1840_inst_ack_1 : boolean;
  signal SLT_f32_u1_1890_inst_req_1 : boolean;
  signal if_stmt_1842_branch_req_0 : boolean;
  signal ADD_f32_f32_1884_inst_ack_0 : boolean;
  signal if_stmt_1842_branch_ack_1 : boolean;
  signal if_stmt_1842_branch_ack_0 : boolean;
  signal type_cast_1954_inst_req_1 : boolean;
  signal type_cast_1954_inst_ack_1 : boolean;
  signal ADD_f32_f32_1884_inst_req_0 : boolean;
  signal SLT_f32_u1_1890_inst_ack_0 : boolean;
  signal SLT_f32_u1_1890_inst_req_0 : boolean;
  signal SGT_f64_u1_1853_inst_req_0 : boolean;
  signal SGT_f64_u1_1853_inst_ack_0 : boolean;
  signal SGT_f64_u1_1853_inst_req_1 : boolean;
  signal SGT_f64_u1_1853_inst_ack_1 : boolean;
  signal ADD_f32_f32_1884_inst_ack_1 : boolean;
  signal ADD_f32_f32_1884_inst_req_1 : boolean;
  signal if_stmt_1855_branch_req_0 : boolean;
  signal if_stmt_1855_branch_ack_1 : boolean;
  signal SUB_u32_u32_2322_inst_req_0 : boolean;
  signal if_stmt_1855_branch_ack_0 : boolean;
  signal ADD_u32_u32_2317_inst_req_1 : boolean;
  signal MUL_f32_f32_1879_inst_req_0 : boolean;
  signal MUL_f32_f32_1879_inst_ack_0 : boolean;
  signal MUL_f32_f32_1879_inst_req_1 : boolean;
  signal MUL_f32_f32_1879_inst_ack_1 : boolean;
  signal AND_u32_u32_2003_inst_req_0 : boolean;
  signal AND_u32_u32_2003_inst_ack_0 : boolean;
  signal AND_u32_u32_2003_inst_req_1 : boolean;
  signal AND_u32_u32_2003_inst_ack_1 : boolean;
  signal OR_u32_u32_2009_inst_req_0 : boolean;
  signal OR_u32_u32_2009_inst_ack_0 : boolean;
  signal OR_u32_u32_2009_inst_req_1 : boolean;
  signal OR_u32_u32_2009_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2015_inst_req_0 : boolean;
  signal LSHR_u32_u32_2015_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2015_inst_req_1 : boolean;
  signal LSHR_u32_u32_2015_inst_ack_1 : boolean;
  signal AND_u32_u32_2021_inst_req_0 : boolean;
  signal AND_u32_u32_2021_inst_ack_0 : boolean;
  signal AND_u32_u32_2021_inst_req_1 : boolean;
  signal AND_u32_u32_2021_inst_ack_1 : boolean;
  signal OR_u32_u32_2027_inst_req_0 : boolean;
  signal OR_u32_u32_2027_inst_ack_0 : boolean;
  signal OR_u32_u32_2027_inst_req_1 : boolean;
  signal OR_u32_u32_2027_inst_ack_1 : boolean;
  signal XOR_u32_u32_2032_inst_req_0 : boolean;
  signal XOR_u32_u32_2032_inst_ack_0 : boolean;
  signal XOR_u32_u32_2032_inst_req_1 : boolean;
  signal XOR_u32_u32_2032_inst_ack_1 : boolean;
  signal AND_u32_u32_2038_inst_req_0 : boolean;
  signal AND_u32_u32_2038_inst_ack_0 : boolean;
  signal AND_u32_u32_2038_inst_req_1 : boolean;
  signal AND_u32_u32_2038_inst_ack_1 : boolean;
  signal if_stmt_2286_branch_ack_1 : boolean;
  signal XOR_u32_u32_2312_inst_ack_0 : boolean;
  signal XOR_u32_u32_2312_inst_req_0 : boolean;
  signal SUB_u32_u32_2043_inst_req_0 : boolean;
  signal SUB_u32_u32_2043_inst_ack_0 : boolean;
  signal SUB_u32_u32_2043_inst_req_1 : boolean;
  signal SUB_u32_u32_2043_inst_ack_1 : boolean;
  signal ADD_u32_u32_2284_inst_ack_1 : boolean;
  signal switch_stmt_2045_branch_default_req_0 : boolean;
  signal switch_stmt_2045_select_expr_0_req_0 : boolean;
  signal switch_stmt_2045_select_expr_0_ack_0 : boolean;
  signal switch_stmt_2045_select_expr_0_req_1 : boolean;
  signal switch_stmt_2045_select_expr_0_ack_1 : boolean;
  signal switch_stmt_2045_branch_0_req_0 : boolean;
  signal OR_u32_u32_2306_inst_ack_1 : boolean;
  signal switch_stmt_2045_select_expr_1_req_0 : boolean;
  signal switch_stmt_2045_select_expr_1_ack_0 : boolean;
  signal OR_u32_u32_2306_inst_req_1 : boolean;
  signal switch_stmt_2045_select_expr_1_req_1 : boolean;
  signal switch_stmt_2045_select_expr_1_ack_1 : boolean;
  signal switch_stmt_2045_branch_1_req_0 : boolean;
  signal AND_u32_u32_2974_inst_ack_1 : boolean;
  signal ADD_u32_u32_2284_inst_req_1 : boolean;
  signal switch_stmt_2045_branch_0_ack_1 : boolean;
  signal switch_stmt_2045_branch_1_ack_1 : boolean;
  signal ADD_u32_u32_2284_inst_ack_0 : boolean;
  signal OR_u32_u32_2306_inst_ack_0 : boolean;
  signal switch_stmt_2045_branch_default_ack_0 : boolean;
  signal ADD_u32_u32_2317_inst_ack_0 : boolean;
  signal OR_u32_u32_2306_inst_req_0 : boolean;
  signal LSHR_u32_u32_2076_inst_req_0 : boolean;
  signal LSHR_u32_u32_2076_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2076_inst_req_1 : boolean;
  signal LSHR_u32_u32_2076_inst_ack_1 : boolean;
  signal ADD_u32_u32_2317_inst_ack_1 : boolean;
  signal AND_u32_u32_2650_inst_req_1 : boolean;
  signal UGT_u32_u1_2081_inst_req_0 : boolean;
  signal UGT_u32_u1_2081_inst_ack_0 : boolean;
  signal UGT_u32_u1_2081_inst_req_1 : boolean;
  signal UGT_u32_u1_2081_inst_ack_1 : boolean;
  signal type_cast_2660_inst_req_0 : boolean;
  signal EQ_u32_u1_2656_inst_req_1 : boolean;
  signal type_cast_2660_inst_req_1 : boolean;
  signal ADD_u32_u32_2284_inst_req_0 : boolean;
  signal if_stmt_2083_branch_req_0 : boolean;
  signal if_stmt_2083_branch_ack_1 : boolean;
  signal if_stmt_2083_branch_ack_0 : boolean;
  signal ADD_u32_u32_2317_inst_req_0 : boolean;
  signal if_stmt_2286_branch_req_0 : boolean;
  signal SHL_u32_u32_2110_inst_req_0 : boolean;
  signal SHL_u32_u32_2110_inst_ack_0 : boolean;
  signal if_stmt_2286_branch_ack_0 : boolean;
  signal SHL_u32_u32_2110_inst_req_1 : boolean;
  signal SHL_u32_u32_2110_inst_ack_1 : boolean;
  signal AND_u32_u32_2650_inst_ack_1 : boolean;
  signal SHL_u32_u32_2116_inst_req_0 : boolean;
  signal SHL_u32_u32_2116_inst_ack_0 : boolean;
  signal SHL_u32_u32_2116_inst_req_1 : boolean;
  signal SHL_u32_u32_2116_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2664_inst_ack_0 : boolean;
  signal ULT_u32_u1_2121_inst_req_0 : boolean;
  signal ULT_u32_u1_2121_inst_ack_0 : boolean;
  signal ULT_u32_u1_2121_inst_req_1 : boolean;
  signal ULT_u32_u1_2121_inst_ack_1 : boolean;
  signal if_stmt_2123_branch_req_0 : boolean;
  signal AND_u32_u32_2650_inst_req_0 : boolean;
  signal if_stmt_2123_branch_ack_1 : boolean;
  signal if_stmt_2123_branch_ack_0 : boolean;
  signal AND_u32_u32_2650_inst_ack_0 : boolean;
  signal EQ_u32_u1_2656_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2664_inst_req_0 : boolean;
  signal type_cast_2660_inst_ack_0 : boolean;
  signal ADD_u32_u32_2158_inst_req_0 : boolean;
  signal ADD_u32_u32_2158_inst_ack_0 : boolean;
  signal ADD_u32_u32_2158_inst_req_1 : boolean;
  signal ADD_u32_u32_2158_inst_ack_1 : boolean;
  signal SUB_u32_u32_2163_inst_req_0 : boolean;
  signal SUB_u32_u32_2163_inst_ack_0 : boolean;
  signal SUB_u32_u32_2163_inst_req_1 : boolean;
  signal SUB_u32_u32_2163_inst_ack_1 : boolean;
  signal type_cast_2660_inst_ack_1 : boolean;
  signal EQ_u32_u1_2656_inst_req_0 : boolean;
  signal ULT_u32_u1_2168_inst_req_0 : boolean;
  signal ULT_u32_u1_2168_inst_ack_0 : boolean;
  signal ULT_u32_u1_2168_inst_req_1 : boolean;
  signal ULT_u32_u1_2168_inst_ack_1 : boolean;
  signal EQ_u32_u1_2656_inst_ack_1 : boolean;
  signal if_stmt_2170_branch_req_0 : boolean;
  signal NEQ_i32_u1_2664_inst_req_1 : boolean;
  signal if_stmt_2170_branch_ack_1 : boolean;
  signal NEQ_i32_u1_2664_inst_ack_1 : boolean;
  signal if_stmt_2170_branch_ack_0 : boolean;
  signal AND_u32_u32_2205_inst_req_0 : boolean;
  signal AND_u32_u32_2205_inst_ack_0 : boolean;
  signal AND_u32_u32_2205_inst_req_1 : boolean;
  signal AND_u32_u32_2205_inst_ack_1 : boolean;
  signal EQ_u32_u1_2211_inst_req_0 : boolean;
  signal EQ_u32_u1_2211_inst_ack_0 : boolean;
  signal EQ_u32_u1_2211_inst_req_1 : boolean;
  signal EQ_u32_u1_2211_inst_ack_1 : boolean;
  signal type_cast_2215_inst_req_0 : boolean;
  signal type_cast_2215_inst_ack_0 : boolean;
  signal type_cast_2215_inst_req_1 : boolean;
  signal type_cast_2215_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2219_inst_req_0 : boolean;
  signal NEQ_i32_u1_2219_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2219_inst_req_1 : boolean;
  signal NEQ_i32_u1_2219_inst_ack_1 : boolean;
  signal AND_u1_u1_2224_inst_req_0 : boolean;
  signal AND_u1_u1_2224_inst_ack_0 : boolean;
  signal AND_u1_u1_2224_inst_req_1 : boolean;
  signal AND_u1_u1_2224_inst_ack_1 : boolean;
  signal if_stmt_2226_branch_req_0 : boolean;
  signal if_stmt_2226_branch_ack_1 : boolean;
  signal if_stmt_2226_branch_ack_0 : boolean;
  signal SHL_u32_u32_2253_inst_req_0 : boolean;
  signal SHL_u32_u32_2253_inst_ack_0 : boolean;
  signal SHL_u32_u32_2253_inst_req_1 : boolean;
  signal SHL_u32_u32_2253_inst_ack_1 : boolean;
  signal AND_u32_u32_2259_inst_req_0 : boolean;
  signal AND_u32_u32_2259_inst_ack_0 : boolean;
  signal AND_u32_u32_2259_inst_req_1 : boolean;
  signal AND_u32_u32_2259_inst_ack_1 : boolean;
  signal EQ_u32_u1_2265_inst_req_0 : boolean;
  signal EQ_u32_u1_2265_inst_ack_0 : boolean;
  signal EQ_u32_u1_2265_inst_req_1 : boolean;
  signal EQ_u32_u1_2265_inst_ack_1 : boolean;
  signal type_cast_2269_inst_req_0 : boolean;
  signal type_cast_2269_inst_ack_0 : boolean;
  signal type_cast_2269_inst_req_1 : boolean;
  signal type_cast_2269_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2273_inst_req_0 : boolean;
  signal NEQ_i32_u1_2273_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2273_inst_req_1 : boolean;
  signal NEQ_i32_u1_2273_inst_ack_1 : boolean;
  signal AND_u1_u1_2278_inst_req_0 : boolean;
  signal AND_u1_u1_2278_inst_ack_0 : boolean;
  signal AND_u1_u1_2278_inst_req_1 : boolean;
  signal AND_u1_u1_2278_inst_ack_1 : boolean;
  signal SUB_u32_u32_2322_inst_req_1 : boolean;
  signal SUB_u32_u32_2322_inst_ack_1 : boolean;
  signal AND_u32_u32_2343_inst_req_0 : boolean;
  signal AND_u32_u32_2343_inst_ack_0 : boolean;
  signal AND_u32_u32_2343_inst_req_1 : boolean;
  signal AND_u32_u32_2343_inst_ack_1 : boolean;
  signal SHL_u32_u32_2349_inst_req_0 : boolean;
  signal SHL_u32_u32_2349_inst_ack_0 : boolean;
  signal SHL_u32_u32_2349_inst_req_1 : boolean;
  signal SHL_u32_u32_2349_inst_ack_1 : boolean;
  signal ADD_u32_u32_2355_inst_req_0 : boolean;
  signal ADD_u32_u32_2355_inst_ack_0 : boolean;
  signal ADD_u32_u32_2355_inst_req_1 : boolean;
  signal ADD_u32_u32_2355_inst_ack_1 : boolean;
  signal OR_u32_u32_2360_inst_req_0 : boolean;
  signal OR_u32_u32_2360_inst_ack_0 : boolean;
  signal OR_u32_u32_2360_inst_req_1 : boolean;
  signal OR_u32_u32_2360_inst_ack_1 : boolean;
  signal OR_u32_u32_2365_inst_req_0 : boolean;
  signal OR_u32_u32_2365_inst_ack_0 : boolean;
  signal OR_u32_u32_2365_inst_req_1 : boolean;
  signal OR_u32_u32_2365_inst_ack_1 : boolean;
  signal type_cast_2369_inst_req_0 : boolean;
  signal type_cast_2369_inst_ack_0 : boolean;
  signal type_cast_2369_inst_req_1 : boolean;
  signal type_cast_2369_inst_ack_1 : boolean;
  signal ADD_f32_f32_2384_inst_req_0 : boolean;
  signal ADD_f32_f32_2384_inst_ack_0 : boolean;
  signal ADD_f32_f32_2384_inst_req_1 : boolean;
  signal ADD_f32_f32_2384_inst_ack_1 : boolean;
  signal MUL_f32_f32_2390_inst_req_0 : boolean;
  signal MUL_f32_f32_2390_inst_ack_0 : boolean;
  signal MUL_f32_f32_2390_inst_req_1 : boolean;
  signal MUL_f32_f32_2390_inst_ack_1 : boolean;
  signal ADD_f32_f32_2395_inst_req_0 : boolean;
  signal ADD_f32_f32_2395_inst_ack_0 : boolean;
  signal ADD_f32_f32_2395_inst_req_1 : boolean;
  signal ADD_f32_f32_2395_inst_ack_1 : boolean;
  signal type_cast_2399_inst_req_0 : boolean;
  signal type_cast_2399_inst_ack_0 : boolean;
  signal type_cast_2399_inst_req_1 : boolean;
  signal type_cast_2399_inst_ack_1 : boolean;
  signal EQ_f32_u1_2405_inst_req_0 : boolean;
  signal EQ_f32_u1_2405_inst_ack_0 : boolean;
  signal EQ_f32_u1_2405_inst_req_1 : boolean;
  signal EQ_f32_u1_2405_inst_ack_1 : boolean;
  signal if_stmt_2407_branch_req_0 : boolean;
  signal if_stmt_2407_branch_ack_1 : boolean;
  signal if_stmt_2407_branch_ack_0 : boolean;
  signal LSHR_u32_u32_2418_inst_req_0 : boolean;
  signal LSHR_u32_u32_2418_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2418_inst_req_1 : boolean;
  signal LSHR_u32_u32_2418_inst_ack_1 : boolean;
  signal AND_u32_u32_2424_inst_req_0 : boolean;
  signal AND_u32_u32_2424_inst_ack_0 : boolean;
  signal AND_u32_u32_2424_inst_req_1 : boolean;
  signal AND_u32_u32_2424_inst_ack_1 : boolean;
  signal LSHR_u32_u32_3002_inst_req_0 : boolean;
  signal LSHR_u32_u32_3002_inst_ack_0 : boolean;
  signal OR_u32_u32_2980_inst_req_1 : boolean;
  signal LSHR_u32_u32_2430_inst_req_0 : boolean;
  signal LSHR_u32_u32_2430_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2430_inst_req_1 : boolean;
  signal LSHR_u32_u32_2430_inst_ack_1 : boolean;
  signal AND_u32_u32_2436_inst_req_0 : boolean;
  signal AND_u32_u32_2436_inst_ack_0 : boolean;
  signal SHL_u32_u32_2968_inst_req_0 : boolean;
  signal AND_u32_u32_2436_inst_req_1 : boolean;
  signal AND_u32_u32_2436_inst_ack_1 : boolean;
  signal SHL_u32_u32_2968_inst_ack_0 : boolean;
  signal SHL_u32_u32_2442_inst_req_0 : boolean;
  signal SHL_u32_u32_2442_inst_ack_0 : boolean;
  signal SHL_u32_u32_2442_inst_req_1 : boolean;
  signal SHL_u32_u32_2442_inst_ack_1 : boolean;
  signal OR_u32_u32_2980_inst_ack_1 : boolean;
  signal type_cast_2962_inst_req_0 : boolean;
  signal AND_u32_u32_2448_inst_req_0 : boolean;
  signal AND_u32_u32_2448_inst_ack_0 : boolean;
  signal type_cast_2962_inst_ack_0 : boolean;
  signal AND_u32_u32_2448_inst_req_1 : boolean;
  signal AND_u32_u32_2448_inst_ack_1 : boolean;
  signal OR_u32_u32_2454_inst_req_0 : boolean;
  signal OR_u32_u32_2454_inst_ack_0 : boolean;
  signal OR_u32_u32_2454_inst_req_1 : boolean;
  signal OR_u32_u32_2454_inst_ack_1 : boolean;
  signal LSHR_u32_u32_2460_inst_req_0 : boolean;
  signal LSHR_u32_u32_2460_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2460_inst_req_1 : boolean;
  signal LSHR_u32_u32_2460_inst_ack_1 : boolean;
  signal OR_u32_u32_2980_inst_ack_0 : boolean;
  signal type_cast_2962_inst_ack_1 : boolean;
  signal SHL_u32_u32_2968_inst_req_1 : boolean;
  signal AND_u32_u32_2974_inst_req_1 : boolean;
  signal SHL_u32_u32_2968_inst_ack_1 : boolean;
  signal AND_u32_u32_2466_inst_req_0 : boolean;
  signal AND_u32_u32_2466_inst_ack_0 : boolean;
  signal AND_u32_u32_2466_inst_req_1 : boolean;
  signal AND_u32_u32_2466_inst_ack_1 : boolean;
  signal OR_u32_u32_2472_inst_req_0 : boolean;
  signal OR_u32_u32_2472_inst_ack_0 : boolean;
  signal OR_u32_u32_2472_inst_req_1 : boolean;
  signal OR_u32_u32_2472_inst_ack_1 : boolean;
  signal XOR_u32_u32_2477_inst_req_0 : boolean;
  signal XOR_u32_u32_2477_inst_ack_0 : boolean;
  signal XOR_u32_u32_2477_inst_req_1 : boolean;
  signal XOR_u32_u32_2477_inst_ack_1 : boolean;
  signal AND_u32_u32_2483_inst_req_0 : boolean;
  signal AND_u32_u32_2483_inst_ack_0 : boolean;
  signal AND_u32_u32_2483_inst_req_1 : boolean;
  signal AND_u32_u32_2483_inst_ack_1 : boolean;
  signal OR_u32_u32_2980_inst_req_0 : boolean;
  signal type_cast_2962_inst_req_1 : boolean;
  signal SUB_u32_u32_2488_inst_req_0 : boolean;
  signal SUB_u32_u32_2488_inst_ack_0 : boolean;
  signal SUB_u32_u32_2488_inst_req_1 : boolean;
  signal SUB_u32_u32_2488_inst_ack_1 : boolean;
  signal switch_stmt_2490_branch_default_req_0 : boolean;
  signal switch_stmt_2490_select_expr_0_req_0 : boolean;
  signal switch_stmt_2490_select_expr_0_ack_0 : boolean;
  signal switch_stmt_2490_select_expr_0_req_1 : boolean;
  signal switch_stmt_2490_select_expr_0_ack_1 : boolean;
  signal switch_stmt_2490_branch_0_req_0 : boolean;
  signal AND_u32_u32_2974_inst_req_0 : boolean;
  signal AND_u32_u32_2974_inst_ack_0 : boolean;
  signal switch_stmt_2490_select_expr_1_req_0 : boolean;
  signal switch_stmt_2490_select_expr_1_ack_0 : boolean;
  signal switch_stmt_2490_select_expr_1_req_1 : boolean;
  signal switch_stmt_2490_select_expr_1_ack_1 : boolean;
  signal switch_stmt_2490_branch_1_req_0 : boolean;
  signal switch_stmt_2490_branch_0_ack_1 : boolean;
  signal switch_stmt_2490_branch_1_ack_1 : boolean;
  signal switch_stmt_2490_branch_default_ack_0 : boolean;
  signal LSHR_u32_u32_2521_inst_req_0 : boolean;
  signal LSHR_u32_u32_2521_inst_ack_0 : boolean;
  signal LSHR_u32_u32_2521_inst_req_1 : boolean;
  signal LSHR_u32_u32_2521_inst_ack_1 : boolean;
  signal UGT_u32_u1_2526_inst_req_0 : boolean;
  signal UGT_u32_u1_2526_inst_ack_0 : boolean;
  signal UGT_u32_u1_2526_inst_req_1 : boolean;
  signal UGT_u32_u1_2526_inst_ack_1 : boolean;
  signal if_stmt_2528_branch_req_0 : boolean;
  signal if_stmt_2528_branch_ack_1 : boolean;
  signal if_stmt_2528_branch_ack_0 : boolean;
  signal SHL_u32_u32_2555_inst_req_0 : boolean;
  signal SHL_u32_u32_2555_inst_ack_0 : boolean;
  signal SHL_u32_u32_2555_inst_req_1 : boolean;
  signal SHL_u32_u32_2555_inst_ack_1 : boolean;
  signal SHL_u32_u32_2561_inst_req_0 : boolean;
  signal SHL_u32_u32_2561_inst_ack_0 : boolean;
  signal SHL_u32_u32_2561_inst_req_1 : boolean;
  signal SHL_u32_u32_2561_inst_ack_1 : boolean;
  signal ULT_u32_u1_2566_inst_req_0 : boolean;
  signal ULT_u32_u1_2566_inst_ack_0 : boolean;
  signal ULT_u32_u1_2566_inst_req_1 : boolean;
  signal ULT_u32_u1_2566_inst_ack_1 : boolean;
  signal if_stmt_2568_branch_req_0 : boolean;
  signal if_stmt_2568_branch_ack_1 : boolean;
  signal if_stmt_2568_branch_ack_0 : boolean;
  signal ADD_u32_u32_2603_inst_req_0 : boolean;
  signal ADD_u32_u32_2603_inst_ack_0 : boolean;
  signal ADD_u32_u32_2603_inst_req_1 : boolean;
  signal ADD_u32_u32_2603_inst_ack_1 : boolean;
  signal SUB_u32_u32_2608_inst_req_0 : boolean;
  signal SUB_u32_u32_2608_inst_ack_0 : boolean;
  signal SUB_u32_u32_2608_inst_req_1 : boolean;
  signal SUB_u32_u32_2608_inst_ack_1 : boolean;
  signal ULT_u32_u1_2613_inst_req_0 : boolean;
  signal ULT_u32_u1_2613_inst_ack_0 : boolean;
  signal ULT_u32_u1_2613_inst_req_1 : boolean;
  signal ULT_u32_u1_2613_inst_ack_1 : boolean;
  signal if_stmt_2615_branch_req_0 : boolean;
  signal if_stmt_2615_branch_ack_1 : boolean;
  signal if_stmt_2615_branch_ack_0 : boolean;
  signal AND_u1_u1_2669_inst_req_0 : boolean;
  signal AND_u1_u1_2669_inst_ack_0 : boolean;
  signal AND_u1_u1_2669_inst_req_1 : boolean;
  signal AND_u1_u1_2669_inst_ack_1 : boolean;
  signal if_stmt_2671_branch_req_0 : boolean;
  signal if_stmt_2671_branch_ack_1 : boolean;
  signal if_stmt_2671_branch_ack_0 : boolean;
  signal SHL_u32_u32_2698_inst_req_0 : boolean;
  signal SHL_u32_u32_2698_inst_ack_0 : boolean;
  signal SHL_u32_u32_2698_inst_req_1 : boolean;
  signal SHL_u32_u32_2698_inst_ack_1 : boolean;
  signal AND_u32_u32_2704_inst_req_0 : boolean;
  signal AND_u32_u32_2704_inst_ack_0 : boolean;
  signal AND_u32_u32_2704_inst_req_1 : boolean;
  signal AND_u32_u32_2704_inst_ack_1 : boolean;
  signal EQ_u32_u1_2710_inst_req_0 : boolean;
  signal EQ_u32_u1_2710_inst_ack_0 : boolean;
  signal EQ_u32_u1_2710_inst_req_1 : boolean;
  signal EQ_u32_u1_2710_inst_ack_1 : boolean;
  signal type_cast_2714_inst_req_0 : boolean;
  signal type_cast_2714_inst_ack_0 : boolean;
  signal type_cast_2714_inst_req_1 : boolean;
  signal type_cast_2714_inst_ack_1 : boolean;
  signal NEQ_i32_u1_2718_inst_req_0 : boolean;
  signal NEQ_i32_u1_2718_inst_ack_0 : boolean;
  signal NEQ_i32_u1_2718_inst_req_1 : boolean;
  signal NEQ_i32_u1_2718_inst_ack_1 : boolean;
  signal AND_u1_u1_2723_inst_req_0 : boolean;
  signal AND_u1_u1_2723_inst_ack_0 : boolean;
  signal AND_u1_u1_2723_inst_req_1 : boolean;
  signal AND_u1_u1_2723_inst_ack_1 : boolean;
  signal ADD_u32_u32_2729_inst_req_0 : boolean;
  signal ADD_u32_u32_2729_inst_ack_0 : boolean;
  signal ADD_u32_u32_2729_inst_req_1 : boolean;
  signal ADD_u32_u32_2729_inst_ack_1 : boolean;
  signal if_stmt_2731_branch_req_0 : boolean;
  signal if_stmt_2731_branch_ack_1 : boolean;
  signal if_stmt_2731_branch_ack_0 : boolean;
  signal OR_u32_u32_2751_inst_req_0 : boolean;
  signal OR_u32_u32_2751_inst_ack_0 : boolean;
  signal OR_u32_u32_2751_inst_req_1 : boolean;
  signal OR_u32_u32_2751_inst_ack_1 : boolean;
  signal XOR_u32_u32_2757_inst_req_0 : boolean;
  signal XOR_u32_u32_2757_inst_ack_0 : boolean;
  signal XOR_u32_u32_2757_inst_req_1 : boolean;
  signal XOR_u32_u32_2757_inst_ack_1 : boolean;
  signal ADD_u32_u32_2762_inst_req_0 : boolean;
  signal ADD_u32_u32_2762_inst_ack_0 : boolean;
  signal ADD_u32_u32_2762_inst_req_1 : boolean;
  signal ADD_u32_u32_2762_inst_ack_1 : boolean;
  signal SUB_u32_u32_2767_inst_req_0 : boolean;
  signal SUB_u32_u32_2767_inst_ack_0 : boolean;
  signal SUB_u32_u32_2767_inst_req_1 : boolean;
  signal SUB_u32_u32_2767_inst_ack_1 : boolean;
  signal AND_u32_u32_2788_inst_req_0 : boolean;
  signal AND_u32_u32_2788_inst_ack_0 : boolean;
  signal AND_u32_u32_2788_inst_req_1 : boolean;
  signal AND_u32_u32_2788_inst_ack_1 : boolean;
  signal SHL_u32_u32_2794_inst_req_0 : boolean;
  signal SHL_u32_u32_2794_inst_ack_0 : boolean;
  signal SHL_u32_u32_2794_inst_req_1 : boolean;
  signal SHL_u32_u32_2794_inst_ack_1 : boolean;
  signal WPIPE_out_data_3311_inst_ack_0 : boolean;
  signal type_cast_3293_inst_req_1 : boolean;
  signal ADD_u32_u32_2800_inst_req_0 : boolean;
  signal ADD_u32_u32_2800_inst_ack_0 : boolean;
  signal type_cast_3293_inst_ack_1 : boolean;
  signal ADD_u32_u32_2800_inst_req_1 : boolean;
  signal ADD_u32_u32_2800_inst_ack_1 : boolean;
  signal MUL_f32_f32_3321_inst_req_0 : boolean;
  signal MUL_f32_f32_3321_inst_ack_0 : boolean;
  signal OR_u32_u32_2805_inst_req_0 : boolean;
  signal OR_u32_u32_2805_inst_ack_0 : boolean;
  signal OR_u32_u32_2805_inst_req_1 : boolean;
  signal OR_u32_u32_2805_inst_ack_1 : boolean;
  signal type_cast_3293_inst_req_0 : boolean;
  signal type_cast_3293_inst_ack_0 : boolean;
  signal OR_u32_u32_2810_inst_req_0 : boolean;
  signal OR_u32_u32_2810_inst_ack_0 : boolean;
  signal OR_u32_u32_2810_inst_req_1 : boolean;
  signal OR_u32_u32_2810_inst_ack_1 : boolean;
  signal WPIPE_out_data_3314_inst_req_0 : boolean;
  signal WPIPE_out_data_3308_inst_req_0 : boolean;
  signal type_cast_2814_inst_req_0 : boolean;
  signal type_cast_2814_inst_ack_0 : boolean;
  signal type_cast_2814_inst_req_1 : boolean;
  signal type_cast_2814_inst_ack_1 : boolean;
  signal WPIPE_out_data_3311_inst_req_0 : boolean;
  signal MUL_f32_f32_2830_inst_req_0 : boolean;
  signal MUL_f32_f32_2830_inst_ack_0 : boolean;
  signal MUL_f32_f32_2830_inst_req_1 : boolean;
  signal MUL_f32_f32_2830_inst_ack_1 : boolean;
  signal WPIPE_out_data_3311_inst_req_1 : boolean;
  signal ADD_f32_f32_2835_inst_req_0 : boolean;
  signal ADD_f32_f32_2835_inst_ack_0 : boolean;
  signal ADD_f32_f32_2835_inst_req_1 : boolean;
  signal ADD_f32_f32_2835_inst_ack_1 : boolean;
  signal WPIPE_out_data_3314_inst_ack_0 : boolean;
  signal WPIPE_out_data_3308_inst_ack_0 : boolean;
  signal SUB_f32_f32_2841_inst_req_0 : boolean;
  signal SUB_f32_f32_2841_inst_ack_0 : boolean;
  signal SUB_f32_f32_2841_inst_req_1 : boolean;
  signal SUB_f32_f32_2841_inst_ack_1 : boolean;
  signal WPIPE_out_data_3308_inst_req_1 : boolean;
  signal WPIPE_out_data_3308_inst_ack_1 : boolean;
  signal MUL_f32_f32_2847_inst_req_0 : boolean;
  signal MUL_f32_f32_2847_inst_ack_0 : boolean;
  signal MUL_f32_f32_2847_inst_req_1 : boolean;
  signal MUL_f32_f32_2847_inst_ack_1 : boolean;
  signal WPIPE_out_data_3311_inst_ack_1 : boolean;
  signal ADD_f32_f32_2852_inst_req_0 : boolean;
  signal ADD_f32_f32_2852_inst_ack_0 : boolean;
  signal ADD_f32_f32_2852_inst_req_1 : boolean;
  signal ADD_f32_f32_2852_inst_ack_1 : boolean;
  signal MUL_f32_f32_3321_inst_req_1 : boolean;
  signal MUL_f32_f32_2858_inst_req_0 : boolean;
  signal MUL_f32_f32_2858_inst_ack_0 : boolean;
  signal MUL_f32_f32_2858_inst_req_1 : boolean;
  signal MUL_f32_f32_2858_inst_ack_1 : boolean;
  signal SLT_f32_u1_2864_inst_req_0 : boolean;
  signal SLT_f32_u1_2864_inst_ack_0 : boolean;
  signal SLT_f32_u1_2864_inst_req_1 : boolean;
  signal SLT_f32_u1_2864_inst_ack_1 : boolean;
  signal if_stmt_2866_branch_req_0 : boolean;
  signal if_stmt_2866_branch_ack_1 : boolean;
  signal if_stmt_2866_branch_ack_0 : boolean;
  signal SGT_f32_u1_2877_inst_req_0 : boolean;
  signal SGT_f32_u1_2877_inst_ack_0 : boolean;
  signal SGT_f32_u1_2877_inst_req_1 : boolean;
  signal SGT_f32_u1_2877_inst_ack_1 : boolean;
  signal if_stmt_2879_branch_req_0 : boolean;
  signal if_stmt_2879_branch_ack_1 : boolean;
  signal if_stmt_2879_branch_ack_0 : boolean;
  signal MUL_f32_f32_2903_inst_req_0 : boolean;
  signal MUL_f32_f32_2903_inst_ack_0 : boolean;
  signal MUL_f32_f32_2903_inst_req_1 : boolean;
  signal MUL_f32_f32_2903_inst_ack_1 : boolean;
  signal ADD_f32_f32_2908_inst_req_0 : boolean;
  signal ADD_f32_f32_2908_inst_ack_0 : boolean;
  signal ADD_f32_f32_2908_inst_req_1 : boolean;
  signal ADD_f32_f32_2908_inst_ack_1 : boolean;
  signal SLT_f32_u1_2914_inst_req_0 : boolean;
  signal SLT_f32_u1_2914_inst_ack_0 : boolean;
  signal SLT_f32_u1_2914_inst_req_1 : boolean;
  signal SLT_f32_u1_2914_inst_ack_1 : boolean;
  signal if_stmt_2916_branch_req_0 : boolean;
  signal if_stmt_2916_branch_ack_1 : boolean;
  signal if_stmt_2916_branch_ack_0 : boolean;
  signal SGT_f32_u1_2927_inst_req_0 : boolean;
  signal SGT_f32_u1_2927_inst_ack_0 : boolean;
  signal SGT_f32_u1_2927_inst_req_1 : boolean;
  signal SGT_f32_u1_2927_inst_ack_1 : boolean;
  signal if_stmt_2929_branch_req_0 : boolean;
  signal if_stmt_2929_branch_ack_1 : boolean;
  signal if_stmt_2929_branch_ack_0 : boolean;
  signal EQ_f32_u1_2940_inst_req_0 : boolean;
  signal EQ_f32_u1_2940_inst_ack_0 : boolean;
  signal EQ_f32_u1_2940_inst_req_1 : boolean;
  signal EQ_f32_u1_2940_inst_ack_1 : boolean;
  signal if_stmt_2942_branch_req_0 : boolean;
  signal if_stmt_2942_branch_ack_1 : boolean;
  signal if_stmt_2942_branch_ack_0 : boolean;
  signal LSHR_u32_u32_3002_inst_req_1 : boolean;
  signal LSHR_u32_u32_3002_inst_ack_1 : boolean;
  signal UGT_u32_u1_3008_inst_req_0 : boolean;
  signal UGT_u32_u1_3008_inst_ack_0 : boolean;
  signal UGT_u32_u1_3008_inst_req_1 : boolean;
  signal UGT_u32_u1_3008_inst_ack_1 : boolean;
  signal if_stmt_3010_branch_req_0 : boolean;
  signal if_stmt_3010_branch_ack_1 : boolean;
  signal if_stmt_3010_branch_ack_0 : boolean;
  signal SHL_u32_u32_3038_inst_req_0 : boolean;
  signal SHL_u32_u32_3038_inst_ack_0 : boolean;
  signal SHL_u32_u32_3038_inst_req_1 : boolean;
  signal SHL_u32_u32_3038_inst_ack_1 : boolean;
  signal SHL_u32_u32_3044_inst_req_0 : boolean;
  signal SHL_u32_u32_3044_inst_ack_0 : boolean;
  signal SHL_u32_u32_3044_inst_req_1 : boolean;
  signal SHL_u32_u32_3044_inst_ack_1 : boolean;
  signal ULT_u32_u1_3049_inst_req_0 : boolean;
  signal ULT_u32_u1_3049_inst_ack_0 : boolean;
  signal ULT_u32_u1_3049_inst_req_1 : boolean;
  signal ULT_u32_u1_3049_inst_ack_1 : boolean;
  signal if_stmt_3051_branch_req_0 : boolean;
  signal if_stmt_3051_branch_ack_1 : boolean;
  signal if_stmt_3051_branch_ack_0 : boolean;
  signal ADD_u32_u32_3087_inst_req_0 : boolean;
  signal ADD_u32_u32_3087_inst_ack_0 : boolean;
  signal ADD_u32_u32_3087_inst_req_1 : boolean;
  signal ADD_u32_u32_3087_inst_ack_1 : boolean;
  signal SUB_u32_u32_3092_inst_req_0 : boolean;
  signal SUB_u32_u32_3092_inst_ack_0 : boolean;
  signal SUB_u32_u32_3092_inst_req_1 : boolean;
  signal SUB_u32_u32_3092_inst_ack_1 : boolean;
  signal ULT_u32_u1_3098_inst_req_0 : boolean;
  signal ULT_u32_u1_3098_inst_ack_0 : boolean;
  signal ULT_u32_u1_3098_inst_req_1 : boolean;
  signal ULT_u32_u1_3098_inst_ack_1 : boolean;
  signal if_stmt_3100_branch_req_0 : boolean;
  signal if_stmt_3100_branch_ack_1 : boolean;
  signal if_stmt_3100_branch_ack_0 : boolean;
  signal LSHR_u32_u32_3116_inst_req_0 : boolean;
  signal LSHR_u32_u32_3116_inst_ack_0 : boolean;
  signal LSHR_u32_u32_3116_inst_req_1 : boolean;
  signal LSHR_u32_u32_3116_inst_ack_1 : boolean;
  signal AND_u32_u32_3122_inst_req_0 : boolean;
  signal AND_u32_u32_3122_inst_ack_0 : boolean;
  signal AND_u32_u32_3122_inst_req_1 : boolean;
  signal AND_u32_u32_3122_inst_ack_1 : boolean;
  signal AND_u32_u32_3128_inst_req_0 : boolean;
  signal AND_u32_u32_3128_inst_ack_0 : boolean;
  signal AND_u32_u32_3128_inst_req_1 : boolean;
  signal AND_u32_u32_3128_inst_ack_1 : boolean;
  signal ADD_u32_u32_3134_inst_req_0 : boolean;
  signal ADD_u32_u32_3134_inst_ack_0 : boolean;
  signal ADD_u32_u32_3134_inst_req_1 : boolean;
  signal ADD_u32_u32_3134_inst_ack_1 : boolean;
  signal AND_u32_u32_3140_inst_req_0 : boolean;
  signal AND_u32_u32_3140_inst_ack_0 : boolean;
  signal AND_u32_u32_3140_inst_req_1 : boolean;
  signal AND_u32_u32_3140_inst_ack_1 : boolean;
  signal WPIPE_out_data_3305_inst_ack_1 : boolean;
  signal WPIPE_out_data_3314_inst_ack_1 : boolean;
  signal WPIPE_out_data_3305_inst_req_1 : boolean;
  signal EQ_u32_u1_3146_inst_req_0 : boolean;
  signal EQ_u32_u1_3146_inst_ack_0 : boolean;
  signal EQ_u32_u1_3146_inst_req_1 : boolean;
  signal EQ_u32_u1_3146_inst_ack_1 : boolean;
  signal WPIPE_out_data_3305_inst_ack_0 : boolean;
  signal WPIPE_out_data_3305_inst_req_0 : boolean;
  signal WPIPE_out_data_3314_inst_req_1 : boolean;
  signal type_cast_3150_inst_req_0 : boolean;
  signal type_cast_3150_inst_ack_0 : boolean;
  signal type_cast_3150_inst_req_1 : boolean;
  signal type_cast_3150_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3154_inst_req_0 : boolean;
  signal NEQ_i32_u1_3154_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3154_inst_req_1 : boolean;
  signal NEQ_i32_u1_3154_inst_ack_1 : boolean;
  signal phi_stmt_2147_req_0 : boolean;
  signal AND_u1_u1_3159_inst_req_0 : boolean;
  signal AND_u1_u1_3159_inst_ack_0 : boolean;
  signal AND_u1_u1_3159_inst_req_1 : boolean;
  signal AND_u1_u1_3159_inst_ack_1 : boolean;
  signal phi_stmt_2184_req_0 : boolean;
  signal if_stmt_3161_branch_req_0 : boolean;
  signal if_stmt_3161_branch_ack_1 : boolean;
  signal if_stmt_3161_branch_ack_0 : boolean;
  signal SHL_u32_u32_3188_inst_req_0 : boolean;
  signal SHL_u32_u32_3188_inst_ack_0 : boolean;
  signal SHL_u32_u32_3188_inst_req_1 : boolean;
  signal SHL_u32_u32_3188_inst_ack_1 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal AND_u32_u32_3194_inst_req_0 : boolean;
  signal AND_u32_u32_3194_inst_ack_0 : boolean;
  signal AND_u32_u32_3194_inst_req_1 : boolean;
  signal AND_u32_u32_3194_inst_ack_1 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal EQ_u32_u1_3200_inst_req_0 : boolean;
  signal EQ_u32_u1_3200_inst_ack_0 : boolean;
  signal EQ_u32_u1_3200_inst_req_1 : boolean;
  signal EQ_u32_u1_3200_inst_ack_1 : boolean;
  signal type_cast_3204_inst_req_0 : boolean;
  signal type_cast_3204_inst_ack_0 : boolean;
  signal type_cast_3204_inst_req_1 : boolean;
  signal type_cast_3204_inst_ack_1 : boolean;
  signal NEQ_i32_u1_3208_inst_req_0 : boolean;
  signal NEQ_i32_u1_3208_inst_ack_0 : boolean;
  signal NEQ_i32_u1_3208_inst_req_1 : boolean;
  signal NEQ_i32_u1_3208_inst_ack_1 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal AND_u1_u1_3213_inst_req_0 : boolean;
  signal AND_u1_u1_3213_inst_ack_0 : boolean;
  signal AND_u1_u1_3213_inst_req_1 : boolean;
  signal AND_u1_u1_3213_inst_ack_1 : boolean;
  signal phi_stmt_2177_req_0 : boolean;
  signal ADD_u32_u32_3219_inst_req_0 : boolean;
  signal ADD_u32_u32_3219_inst_ack_0 : boolean;
  signal ADD_u32_u32_3219_inst_req_1 : boolean;
  signal ADD_u32_u32_3219_inst_ack_1 : boolean;
  signal if_stmt_3221_branch_req_0 : boolean;
  signal if_stmt_3221_branch_ack_1 : boolean;
  signal if_stmt_3221_branch_ack_0 : boolean;
  signal ADD_u32_u32_3241_inst_req_0 : boolean;
  signal ADD_u32_u32_3241_inst_ack_0 : boolean;
  signal ADD_u32_u32_3241_inst_req_1 : boolean;
  signal ADD_u32_u32_3241_inst_ack_1 : boolean;
  signal SUB_u32_u32_3246_inst_req_0 : boolean;
  signal SUB_u32_u32_3246_inst_ack_0 : boolean;
  signal SUB_u32_u32_3246_inst_req_1 : boolean;
  signal SUB_u32_u32_3246_inst_ack_1 : boolean;
  signal AND_u32_u32_3267_inst_req_0 : boolean;
  signal AND_u32_u32_3267_inst_ack_0 : boolean;
  signal AND_u32_u32_3267_inst_req_1 : boolean;
  signal AND_u32_u32_3267_inst_ack_1 : boolean;
  signal SHL_u32_u32_3273_inst_req_0 : boolean;
  signal SHL_u32_u32_3273_inst_ack_0 : boolean;
  signal SHL_u32_u32_3273_inst_req_1 : boolean;
  signal SHL_u32_u32_3273_inst_ack_1 : boolean;
  signal ADD_u32_u32_3279_inst_req_0 : boolean;
  signal ADD_u32_u32_3279_inst_ack_0 : boolean;
  signal ADD_u32_u32_3279_inst_req_1 : boolean;
  signal ADD_u32_u32_3279_inst_ack_1 : boolean;
  signal OR_u32_u32_3284_inst_req_0 : boolean;
  signal OR_u32_u32_3284_inst_ack_0 : boolean;
  signal OR_u32_u32_3284_inst_req_1 : boolean;
  signal OR_u32_u32_3284_inst_ack_1 : boolean;
  signal OR_u32_u32_3289_inst_req_0 : boolean;
  signal OR_u32_u32_3289_inst_ack_0 : boolean;
  signal OR_u32_u32_3289_inst_req_1 : boolean;
  signal OR_u32_u32_3289_inst_ack_1 : boolean;
  signal MUL_f32_f32_3321_inst_ack_1 : boolean;
  signal MUL_f32_f32_3327_inst_req_0 : boolean;
  signal MUL_f32_f32_3327_inst_ack_0 : boolean;
  signal MUL_f32_f32_3327_inst_req_1 : boolean;
  signal MUL_f32_f32_3327_inst_ack_1 : boolean;
  signal MUL_f32_f32_3333_inst_req_0 : boolean;
  signal MUL_f32_f32_3333_inst_ack_0 : boolean;
  signal MUL_f32_f32_3333_inst_req_1 : boolean;
  signal MUL_f32_f32_3333_inst_ack_1 : boolean;
  signal phi_stmt_1697_req_0 : boolean;
  signal phi_stmt_1683_req_0 : boolean;
  signal phi_stmt_1704_req_0 : boolean;
  signal phi_stmt_1676_req_0 : boolean;
  signal phi_stmt_1711_req_0 : boolean;
  signal phi_stmt_1669_req_0 : boolean;
  signal phi_stmt_1690_req_0 : boolean;
  signal phi_stmt_1662_req_0 : boolean;
  signal type_cast_1703_inst_req_0 : boolean;
  signal type_cast_1703_inst_ack_0 : boolean;
  signal type_cast_1703_inst_req_1 : boolean;
  signal type_cast_1703_inst_ack_1 : boolean;
  signal phi_stmt_1697_req_1 : boolean;
  signal type_cast_1689_inst_req_0 : boolean;
  signal type_cast_1689_inst_ack_0 : boolean;
  signal type_cast_1689_inst_req_1 : boolean;
  signal type_cast_1689_inst_ack_1 : boolean;
  signal phi_stmt_1683_req_1 : boolean;
  signal type_cast_1710_inst_req_0 : boolean;
  signal type_cast_1710_inst_ack_0 : boolean;
  signal type_cast_1710_inst_req_1 : boolean;
  signal type_cast_1710_inst_ack_1 : boolean;
  signal phi_stmt_1704_req_1 : boolean;
  signal type_cast_1682_inst_req_0 : boolean;
  signal type_cast_1682_inst_ack_0 : boolean;
  signal type_cast_1682_inst_req_1 : boolean;
  signal type_cast_1682_inst_ack_1 : boolean;
  signal phi_stmt_1676_req_1 : boolean;
  signal type_cast_1717_inst_req_0 : boolean;
  signal type_cast_1717_inst_ack_0 : boolean;
  signal type_cast_1717_inst_req_1 : boolean;
  signal type_cast_1717_inst_ack_1 : boolean;
  signal phi_stmt_1711_req_1 : boolean;
  signal type_cast_1675_inst_req_0 : boolean;
  signal type_cast_1675_inst_ack_0 : boolean;
  signal type_cast_1675_inst_req_1 : boolean;
  signal type_cast_1675_inst_ack_1 : boolean;
  signal phi_stmt_1669_req_1 : boolean;
  signal type_cast_1696_inst_req_0 : boolean;
  signal type_cast_1696_inst_ack_0 : boolean;
  signal type_cast_1696_inst_req_1 : boolean;
  signal type_cast_1696_inst_ack_1 : boolean;
  signal phi_stmt_1690_req_1 : boolean;
  signal type_cast_1668_inst_req_0 : boolean;
  signal type_cast_1668_inst_ack_0 : boolean;
  signal type_cast_1668_inst_req_1 : boolean;
  signal type_cast_1668_inst_ack_1 : boolean;
  signal phi_stmt_1662_req_1 : boolean;
  signal phi_stmt_1662_ack_0 : boolean;
  signal phi_stmt_1669_ack_0 : boolean;
  signal phi_stmt_1676_ack_0 : boolean;
  signal phi_stmt_1683_ack_0 : boolean;
  signal phi_stmt_1690_ack_0 : boolean;
  signal phi_stmt_1697_ack_0 : boolean;
  signal phi_stmt_1704_ack_0 : boolean;
  signal phi_stmt_1711_ack_0 : boolean;
  signal type_cast_1794_inst_req_0 : boolean;
  signal type_cast_1794_inst_ack_0 : boolean;
  signal type_cast_1794_inst_req_1 : boolean;
  signal type_cast_1794_inst_ack_1 : boolean;
  signal phi_stmt_1791_req_0 : boolean;
  signal type_cast_1798_inst_req_0 : boolean;
  signal type_cast_1798_inst_ack_0 : boolean;
  signal type_cast_1798_inst_req_1 : boolean;
  signal type_cast_1798_inst_ack_1 : boolean;
  signal phi_stmt_1791_req_2 : boolean;
  signal type_cast_1796_inst_req_0 : boolean;
  signal type_cast_1796_inst_ack_0 : boolean;
  signal type_cast_1796_inst_req_1 : boolean;
  signal type_cast_1796_inst_ack_1 : boolean;
  signal phi_stmt_1791_req_1 : boolean;
  signal phi_stmt_1791_ack_0 : boolean;
  signal phi_stmt_1864_req_1 : boolean;
  signal phi_stmt_2147_ack_0 : boolean;
  signal phi_stmt_2141_ack_0 : boolean;
  signal phi_stmt_1864_req_2 : boolean;
  signal phi_stmt_2147_req_1 : boolean;
  signal type_cast_2153_inst_ack_1 : boolean;
  signal type_cast_1867_inst_req_0 : boolean;
  signal type_cast_1867_inst_ack_0 : boolean;
  signal type_cast_2153_inst_req_1 : boolean;
  signal type_cast_1867_inst_req_1 : boolean;
  signal type_cast_1867_inst_ack_1 : boolean;
  signal phi_stmt_1864_req_0 : boolean;
  signal phi_stmt_1864_ack_0 : boolean;
  signal type_cast_2153_inst_ack_0 : boolean;
  signal phi_stmt_2141_req_0 : boolean;
  signal type_cast_2153_inst_req_0 : boolean;
  signal type_cast_1923_inst_req_0 : boolean;
  signal type_cast_1923_inst_ack_0 : boolean;
  signal type_cast_1923_inst_req_1 : boolean;
  signal type_cast_1923_inst_ack_1 : boolean;
  signal phi_stmt_1920_req_0 : boolean;
  signal phi_stmt_2141_req_1 : boolean;
  signal type_cast_2146_inst_ack_1 : boolean;
  signal phi_stmt_1920_req_1 : boolean;
  signal type_cast_2146_inst_req_1 : boolean;
  signal type_cast_2146_inst_ack_0 : boolean;
  signal type_cast_2146_inst_req_0 : boolean;
  signal phi_stmt_1920_req_2 : boolean;
  signal phi_stmt_2177_ack_0 : boolean;
  signal phi_stmt_1920_ack_0 : boolean;
  signal phi_stmt_2064_req_1 : boolean;
  signal type_cast_2144_inst_ack_1 : boolean;
  signal type_cast_2063_inst_req_0 : boolean;
  signal type_cast_2063_inst_ack_0 : boolean;
  signal type_cast_2063_inst_req_1 : boolean;
  signal type_cast_2063_inst_ack_1 : boolean;
  signal phi_stmt_2058_req_1 : boolean;
  signal type_cast_2067_inst_req_0 : boolean;
  signal type_cast_2067_inst_ack_0 : boolean;
  signal type_cast_2067_inst_req_1 : boolean;
  signal type_cast_2067_inst_ack_1 : boolean;
  signal type_cast_2774_inst_ack_1 : boolean;
  signal phi_stmt_2064_req_0 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal phi_stmt_2058_req_0 : boolean;
  signal phi_stmt_2058_ack_0 : boolean;
  signal phi_stmt_2064_ack_0 : boolean;
  signal type_cast_2101_inst_req_0 : boolean;
  signal type_cast_2101_inst_ack_0 : boolean;
  signal type_cast_2101_inst_req_1 : boolean;
  signal type_cast_2101_inst_ack_1 : boolean;
  signal phi_stmt_2098_req_0 : boolean;
  signal type_cast_2095_inst_req_0 : boolean;
  signal type_cast_2095_inst_ack_0 : boolean;
  signal type_cast_2095_inst_req_1 : boolean;
  signal type_cast_2095_inst_ack_1 : boolean;
  signal phi_stmt_2092_req_0 : boolean;
  signal phi_stmt_2098_req_1 : boolean;
  signal type_cast_2097_inst_req_0 : boolean;
  signal type_cast_2097_inst_ack_0 : boolean;
  signal type_cast_2097_inst_req_1 : boolean;
  signal type_cast_2097_inst_ack_1 : boolean;
  signal phi_stmt_2092_req_1 : boolean;
  signal phi_stmt_2092_ack_0 : boolean;
  signal phi_stmt_2098_ack_0 : boolean;
  signal type_cast_2133_inst_req_0 : boolean;
  signal type_cast_2133_inst_ack_0 : boolean;
  signal type_cast_2133_inst_req_1 : boolean;
  signal type_cast_2133_inst_ack_1 : boolean;
  signal phi_stmt_2130_req_0 : boolean;
  signal type_cast_2137_inst_req_0 : boolean;
  signal type_cast_2137_inst_ack_0 : boolean;
  signal type_cast_2137_inst_req_1 : boolean;
  signal type_cast_2137_inst_ack_1 : boolean;
  signal phi_stmt_2134_req_0 : boolean;
  signal phi_stmt_2130_ack_0 : boolean;
  signal phi_stmt_2134_ack_0 : boolean;
  signal type_cast_2144_inst_req_0 : boolean;
  signal type_cast_2144_inst_ack_0 : boolean;
  signal type_cast_2144_inst_req_1 : boolean;
  signal type_cast_2190_inst_req_0 : boolean;
  signal type_cast_2190_inst_ack_0 : boolean;
  signal type_cast_2190_inst_req_1 : boolean;
  signal type_cast_2190_inst_ack_1 : boolean;
  signal phi_stmt_2184_req_1 : boolean;
  signal phi_stmt_2184_ack_0 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_1 : boolean;
  signal type_cast_2197_inst_req_0 : boolean;
  signal type_cast_2197_inst_ack_0 : boolean;
  signal type_cast_2197_inst_req_1 : boolean;
  signal type_cast_2197_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_0 : boolean;
  signal phi_stmt_2194_ack_0 : boolean;
  signal type_cast_2238_inst_req_0 : boolean;
  signal type_cast_2238_inst_ack_0 : boolean;
  signal type_cast_2238_inst_req_1 : boolean;
  signal type_cast_2238_inst_ack_1 : boolean;
  signal phi_stmt_2235_req_0 : boolean;
  signal type_cast_2245_inst_req_0 : boolean;
  signal type_cast_2245_inst_ack_0 : boolean;
  signal type_cast_2245_inst_req_1 : boolean;
  signal type_cast_2245_inst_ack_1 : boolean;
  signal phi_stmt_2242_req_0 : boolean;
  signal phi_stmt_2235_req_1 : boolean;
  signal type_cast_2247_inst_req_0 : boolean;
  signal type_cast_2247_inst_ack_0 : boolean;
  signal type_cast_2247_inst_req_1 : boolean;
  signal type_cast_2247_inst_ack_1 : boolean;
  signal phi_stmt_2242_req_1 : boolean;
  signal phi_stmt_2235_ack_0 : boolean;
  signal phi_stmt_2242_ack_0 : boolean;
  signal type_cast_2296_inst_req_0 : boolean;
  signal type_cast_2296_inst_ack_0 : boolean;
  signal type_cast_2296_inst_req_1 : boolean;
  signal type_cast_2296_inst_ack_1 : boolean;
  signal phi_stmt_2293_req_0 : boolean;
  signal type_cast_2300_inst_req_0 : boolean;
  signal type_cast_2300_inst_ack_0 : boolean;
  signal type_cast_2300_inst_req_1 : boolean;
  signal type_cast_2300_inst_ack_1 : boolean;
  signal phi_stmt_2297_req_0 : boolean;
  signal phi_stmt_2293_ack_0 : boolean;
  signal phi_stmt_2297_ack_0 : boolean;
  signal type_cast_2331_inst_req_0 : boolean;
  signal type_cast_2331_inst_ack_0 : boolean;
  signal type_cast_2331_inst_req_1 : boolean;
  signal type_cast_2331_inst_ack_1 : boolean;
  signal phi_stmt_2326_req_1 : boolean;
  signal type_cast_2337_inst_req_0 : boolean;
  signal type_cast_2337_inst_ack_0 : boolean;
  signal type_cast_2337_inst_req_1 : boolean;
  signal type_cast_2337_inst_ack_1 : boolean;
  signal phi_stmt_2332_req_1 : boolean;
  signal type_cast_2329_inst_req_0 : boolean;
  signal type_cast_2329_inst_ack_0 : boolean;
  signal type_cast_2329_inst_req_1 : boolean;
  signal type_cast_2329_inst_ack_1 : boolean;
  signal phi_stmt_2326_req_0 : boolean;
  signal type_cast_2335_inst_req_0 : boolean;
  signal type_cast_2335_inst_ack_0 : boolean;
  signal type_cast_2335_inst_req_1 : boolean;
  signal type_cast_2335_inst_ack_1 : boolean;
  signal phi_stmt_2332_req_0 : boolean;
  signal phi_stmt_2326_ack_0 : boolean;
  signal phi_stmt_2332_ack_0 : boolean;
  signal phi_stmt_2373_req_1 : boolean;
  signal type_cast_2376_inst_req_0 : boolean;
  signal type_cast_2376_inst_ack_0 : boolean;
  signal type_cast_2376_inst_req_1 : boolean;
  signal type_cast_2376_inst_ack_1 : boolean;
  signal phi_stmt_2373_req_0 : boolean;
  signal phi_stmt_2373_ack_0 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_1 : boolean;
  signal phi_stmt_2509_req_1 : boolean;
  signal type_cast_2506_inst_req_0 : boolean;
  signal type_cast_2506_inst_ack_0 : boolean;
  signal type_cast_2506_inst_req_1 : boolean;
  signal type_cast_2506_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_0 : boolean;
  signal type_cast_2512_inst_req_0 : boolean;
  signal type_cast_2512_inst_ack_0 : boolean;
  signal type_cast_2512_inst_req_1 : boolean;
  signal type_cast_2512_inst_ack_1 : boolean;
  signal phi_stmt_2509_req_0 : boolean;
  signal phi_stmt_2503_ack_0 : boolean;
  signal phi_stmt_2509_ack_0 : boolean;
  signal type_cast_2540_inst_req_0 : boolean;
  signal type_cast_2540_inst_ack_0 : boolean;
  signal type_cast_2540_inst_req_1 : boolean;
  signal type_cast_2540_inst_ack_1 : boolean;
  signal phi_stmt_2537_req_0 : boolean;
  signal type_cast_2546_inst_req_0 : boolean;
  signal type_cast_2546_inst_ack_0 : boolean;
  signal type_cast_2546_inst_req_1 : boolean;
  signal type_cast_2546_inst_ack_1 : boolean;
  signal phi_stmt_2543_req_0 : boolean;
  signal type_cast_2542_inst_req_0 : boolean;
  signal type_cast_2542_inst_ack_0 : boolean;
  signal type_cast_2542_inst_req_1 : boolean;
  signal type_cast_2542_inst_ack_1 : boolean;
  signal phi_stmt_2537_req_1 : boolean;
  signal phi_stmt_2543_req_1 : boolean;
  signal phi_stmt_2537_ack_0 : boolean;
  signal phi_stmt_2543_ack_0 : boolean;
  signal type_cast_2578_inst_req_0 : boolean;
  signal type_cast_2578_inst_ack_0 : boolean;
  signal type_cast_2578_inst_req_1 : boolean;
  signal type_cast_2578_inst_ack_1 : boolean;
  signal phi_stmt_2575_req_0 : boolean;
  signal type_cast_2582_inst_req_0 : boolean;
  signal type_cast_2582_inst_ack_0 : boolean;
  signal type_cast_2582_inst_req_1 : boolean;
  signal type_cast_2582_inst_ack_1 : boolean;
  signal phi_stmt_2579_req_0 : boolean;
  signal phi_stmt_2575_ack_0 : boolean;
  signal phi_stmt_2579_ack_0 : boolean;
  signal type_cast_2589_inst_req_0 : boolean;
  signal type_cast_2589_inst_ack_0 : boolean;
  signal type_cast_2589_inst_req_1 : boolean;
  signal type_cast_2589_inst_ack_1 : boolean;
  signal phi_stmt_2586_req_0 : boolean;
  signal phi_stmt_2592_req_0 : boolean;
  signal type_cast_2774_inst_req_1 : boolean;
  signal phi_stmt_2818_ack_0 : boolean;
  signal type_cast_2591_inst_req_0 : boolean;
  signal type_cast_2591_inst_ack_0 : boolean;
  signal type_cast_2591_inst_req_1 : boolean;
  signal type_cast_2591_inst_ack_1 : boolean;
  signal phi_stmt_2586_req_1 : boolean;
  signal phi_stmt_2818_req_0 : boolean;
  signal type_cast_2821_inst_ack_1 : boolean;
  signal type_cast_2598_inst_req_0 : boolean;
  signal type_cast_2598_inst_ack_0 : boolean;
  signal type_cast_2821_inst_req_1 : boolean;
  signal type_cast_2598_inst_req_1 : boolean;
  signal type_cast_2598_inst_ack_1 : boolean;
  signal phi_stmt_2592_req_1 : boolean;
  signal phi_stmt_2586_ack_0 : boolean;
  signal phi_stmt_2592_ack_0 : boolean;
  signal type_cast_2821_inst_ack_0 : boolean;
  signal type_cast_2821_inst_req_0 : boolean;
  signal type_cast_2625_inst_req_0 : boolean;
  signal type_cast_2625_inst_ack_0 : boolean;
  signal type_cast_2625_inst_req_1 : boolean;
  signal type_cast_2625_inst_ack_1 : boolean;
  signal phi_stmt_2622_req_0 : boolean;
  signal type_cast_2774_inst_ack_0 : boolean;
  signal phi_stmt_2622_ack_0 : boolean;
  signal type_cast_2774_inst_req_0 : boolean;
  signal phi_stmt_2818_req_1 : boolean;
  signal phi_stmt_2629_req_0 : boolean;
  signal type_cast_2635_inst_req_0 : boolean;
  signal type_cast_2635_inst_ack_0 : boolean;
  signal type_cast_2635_inst_req_1 : boolean;
  signal type_cast_2635_inst_ack_1 : boolean;
  signal phi_stmt_2629_req_1 : boolean;
  signal phi_stmt_2629_ack_0 : boolean;
  signal type_cast_2644_inst_req_0 : boolean;
  signal type_cast_2644_inst_ack_0 : boolean;
  signal type_cast_2644_inst_req_1 : boolean;
  signal type_cast_2644_inst_ack_1 : boolean;
  signal phi_stmt_2639_req_1 : boolean;
  signal type_cast_2642_inst_req_0 : boolean;
  signal type_cast_2642_inst_ack_0 : boolean;
  signal phi_stmt_2777_ack_0 : boolean;
  signal type_cast_2642_inst_req_1 : boolean;
  signal type_cast_2642_inst_ack_1 : boolean;
  signal phi_stmt_2771_ack_0 : boolean;
  signal phi_stmt_2777_req_0 : boolean;
  signal phi_stmt_2639_req_0 : boolean;
  signal phi_stmt_2639_ack_0 : boolean;
  signal type_cast_2683_inst_req_0 : boolean;
  signal type_cast_2683_inst_ack_0 : boolean;
  signal type_cast_2683_inst_req_1 : boolean;
  signal type_cast_2683_inst_ack_1 : boolean;
  signal phi_stmt_2680_req_0 : boolean;
  signal type_cast_2690_inst_req_0 : boolean;
  signal type_cast_2690_inst_ack_0 : boolean;
  signal type_cast_2780_inst_ack_1 : boolean;
  signal type_cast_2690_inst_req_1 : boolean;
  signal type_cast_2690_inst_ack_1 : boolean;
  signal type_cast_2780_inst_req_1 : boolean;
  signal type_cast_2780_inst_ack_0 : boolean;
  signal phi_stmt_2687_req_0 : boolean;
  signal type_cast_2780_inst_req_0 : boolean;
  signal phi_stmt_2680_req_1 : boolean;
  signal phi_stmt_2771_req_0 : boolean;
  signal type_cast_2692_inst_req_0 : boolean;
  signal type_cast_2692_inst_ack_0 : boolean;
  signal type_cast_2692_inst_req_1 : boolean;
  signal type_cast_2692_inst_ack_1 : boolean;
  signal phi_stmt_2687_req_1 : boolean;
  signal phi_stmt_2680_ack_0 : boolean;
  signal phi_stmt_2687_ack_0 : boolean;
  signal type_cast_2741_inst_req_0 : boolean;
  signal type_cast_2741_inst_ack_0 : boolean;
  signal type_cast_2741_inst_req_1 : boolean;
  signal type_cast_2741_inst_ack_1 : boolean;
  signal phi_stmt_2738_req_0 : boolean;
  signal type_cast_2745_inst_req_0 : boolean;
  signal type_cast_2745_inst_ack_0 : boolean;
  signal type_cast_2745_inst_req_1 : boolean;
  signal type_cast_2745_inst_ack_1 : boolean;
  signal phi_stmt_2742_req_0 : boolean;
  signal phi_stmt_2738_ack_0 : boolean;
  signal phi_stmt_2742_ack_0 : boolean;
  signal type_cast_2776_inst_req_0 : boolean;
  signal type_cast_2776_inst_ack_0 : boolean;
  signal type_cast_2776_inst_req_1 : boolean;
  signal type_cast_2776_inst_ack_1 : boolean;
  signal phi_stmt_2771_req_1 : boolean;
  signal type_cast_2782_inst_req_0 : boolean;
  signal type_cast_2782_inst_ack_0 : boolean;
  signal type_cast_2782_inst_req_1 : boolean;
  signal type_cast_2782_inst_ack_1 : boolean;
  signal phi_stmt_2777_req_1 : boolean;
  signal phi_stmt_2888_req_2 : boolean;
  signal type_cast_2891_inst_req_0 : boolean;
  signal type_cast_2891_inst_ack_0 : boolean;
  signal type_cast_2891_inst_req_1 : boolean;
  signal type_cast_2891_inst_ack_1 : boolean;
  signal phi_stmt_2888_req_0 : boolean;
  signal phi_stmt_2888_req_1 : boolean;
  signal phi_stmt_2888_ack_0 : boolean;
  signal phi_stmt_2949_req_1 : boolean;
  signal phi_stmt_2949_req_2 : boolean;
  signal type_cast_2952_inst_req_0 : boolean;
  signal type_cast_2952_inst_ack_0 : boolean;
  signal type_cast_2952_inst_req_1 : boolean;
  signal type_cast_2952_inst_ack_1 : boolean;
  signal phi_stmt_2949_req_0 : boolean;
  signal phi_stmt_2949_ack_0 : boolean;
  signal type_cast_2987_inst_req_0 : boolean;
  signal type_cast_2987_inst_ack_0 : boolean;
  signal type_cast_2987_inst_req_1 : boolean;
  signal type_cast_2987_inst_ack_1 : boolean;
  signal phi_stmt_2984_req_0 : boolean;
  signal type_cast_2993_inst_req_0 : boolean;
  signal type_cast_2993_inst_ack_0 : boolean;
  signal type_cast_2993_inst_req_1 : boolean;
  signal type_cast_2993_inst_ack_1 : boolean;
  signal phi_stmt_2990_req_0 : boolean;
  signal type_cast_2989_inst_req_0 : boolean;
  signal type_cast_2989_inst_ack_0 : boolean;
  signal type_cast_2989_inst_req_1 : boolean;
  signal type_cast_2989_inst_ack_1 : boolean;
  signal phi_stmt_2984_req_1 : boolean;
  signal phi_stmt_2990_req_1 : boolean;
  signal phi_stmt_2984_ack_0 : boolean;
  signal phi_stmt_2990_ack_0 : boolean;
  signal type_cast_3022_inst_req_0 : boolean;
  signal type_cast_3022_inst_ack_0 : boolean;
  signal type_cast_3022_inst_req_1 : boolean;
  signal type_cast_3022_inst_ack_1 : boolean;
  signal phi_stmt_3019_req_0 : boolean;
  signal type_cast_3029_inst_req_0 : boolean;
  signal type_cast_3029_inst_ack_0 : boolean;
  signal type_cast_3029_inst_req_1 : boolean;
  signal type_cast_3029_inst_ack_1 : boolean;
  signal phi_stmt_3026_req_0 : boolean;
  signal phi_stmt_3019_req_1 : boolean;
  signal phi_stmt_3026_req_1 : boolean;
  signal phi_stmt_3019_ack_0 : boolean;
  signal phi_stmt_3026_ack_0 : boolean;
  signal type_cast_3061_inst_req_0 : boolean;
  signal type_cast_3061_inst_ack_0 : boolean;
  signal type_cast_3061_inst_req_1 : boolean;
  signal type_cast_3061_inst_ack_1 : boolean;
  signal phi_stmt_3058_req_0 : boolean;
  signal type_cast_3065_inst_req_0 : boolean;
  signal type_cast_3065_inst_ack_0 : boolean;
  signal type_cast_3065_inst_req_1 : boolean;
  signal type_cast_3065_inst_ack_1 : boolean;
  signal phi_stmt_3062_req_0 : boolean;
  signal phi_stmt_3058_ack_0 : boolean;
  signal phi_stmt_3062_ack_0 : boolean;
  signal phi_stmt_3069_req_0 : boolean;
  signal phi_stmt_3076_req_0 : boolean;
  signal type_cast_3075_inst_req_0 : boolean;
  signal type_cast_3075_inst_ack_0 : boolean;
  signal type_cast_3075_inst_req_1 : boolean;
  signal type_cast_3075_inst_ack_1 : boolean;
  signal phi_stmt_3069_req_1 : boolean;
  signal type_cast_3082_inst_req_0 : boolean;
  signal type_cast_3082_inst_ack_0 : boolean;
  signal type_cast_3082_inst_req_1 : boolean;
  signal type_cast_3082_inst_ack_1 : boolean;
  signal phi_stmt_3076_req_1 : boolean;
  signal phi_stmt_3069_ack_0 : boolean;
  signal phi_stmt_3076_ack_0 : boolean;
  signal type_cast_3110_inst_req_0 : boolean;
  signal type_cast_3110_inst_ack_0 : boolean;
  signal type_cast_3110_inst_req_1 : boolean;
  signal type_cast_3110_inst_ack_1 : boolean;
  signal phi_stmt_3107_req_0 : boolean;
  signal phi_stmt_3107_ack_0 : boolean;
  signal type_cast_3173_inst_req_0 : boolean;
  signal type_cast_3173_inst_ack_0 : boolean;
  signal type_cast_3173_inst_req_1 : boolean;
  signal type_cast_3173_inst_ack_1 : boolean;
  signal phi_stmt_3170_req_0 : boolean;
  signal type_cast_3180_inst_req_0 : boolean;
  signal type_cast_3180_inst_ack_0 : boolean;
  signal type_cast_3180_inst_req_1 : boolean;
  signal type_cast_3180_inst_ack_1 : boolean;
  signal phi_stmt_3177_req_0 : boolean;
  signal phi_stmt_3170_req_1 : boolean;
  signal type_cast_3182_inst_req_0 : boolean;
  signal type_cast_3182_inst_ack_0 : boolean;
  signal type_cast_3182_inst_req_1 : boolean;
  signal type_cast_3182_inst_ack_1 : boolean;
  signal phi_stmt_3177_req_1 : boolean;
  signal phi_stmt_3170_ack_0 : boolean;
  signal phi_stmt_3177_ack_0 : boolean;
  signal type_cast_3235_inst_req_0 : boolean;
  signal type_cast_3235_inst_ack_0 : boolean;
  signal type_cast_3235_inst_req_1 : boolean;
  signal type_cast_3235_inst_ack_1 : boolean;
  signal phi_stmt_3232_req_0 : boolean;
  signal type_cast_3231_inst_req_0 : boolean;
  signal type_cast_3231_inst_ack_0 : boolean;
  signal type_cast_3231_inst_req_1 : boolean;
  signal type_cast_3231_inst_ack_1 : boolean;
  signal phi_stmt_3228_req_0 : boolean;
  signal phi_stmt_3228_ack_0 : boolean;
  signal phi_stmt_3232_ack_0 : boolean;
  signal type_cast_3255_inst_req_0 : boolean;
  signal type_cast_3255_inst_ack_0 : boolean;
  signal type_cast_3255_inst_req_1 : boolean;
  signal type_cast_3255_inst_ack_1 : boolean;
  signal phi_stmt_3250_req_1 : boolean;
  signal type_cast_3261_inst_req_0 : boolean;
  signal type_cast_3261_inst_ack_0 : boolean;
  signal type_cast_3261_inst_req_1 : boolean;
  signal type_cast_3261_inst_ack_1 : boolean;
  signal phi_stmt_3256_req_1 : boolean;
  signal type_cast_3253_inst_req_0 : boolean;
  signal type_cast_3253_inst_ack_0 : boolean;
  signal type_cast_3253_inst_req_1 : boolean;
  signal type_cast_3253_inst_ack_1 : boolean;
  signal phi_stmt_3250_req_0 : boolean;
  signal type_cast_3259_inst_req_0 : boolean;
  signal type_cast_3259_inst_ack_0 : boolean;
  signal type_cast_3259_inst_req_1 : boolean;
  signal type_cast_3259_inst_ack_1 : boolean;
  signal phi_stmt_3256_req_0 : boolean;
  signal phi_stmt_3250_ack_0 : boolean;
  signal phi_stmt_3256_ack_0 : boolean;
  signal phi_stmt_3297_req_1 : boolean;
  signal type_cast_3300_inst_req_0 : boolean;
  signal type_cast_3300_inst_ack_0 : boolean;
  signal type_cast_3300_inst_req_1 : boolean;
  signal type_cast_3300_inst_ack_1 : boolean;
  signal phi_stmt_3297_req_0 : boolean;
  signal phi_stmt_3297_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "vector_control_daemon_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  vector_control_daemon_CP_8401_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "vector_control_daemon_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0, 
      kill_counter_range => 1) -- 
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      kill => default_zero_sig,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= vector_control_daemon_CP_8401_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= vector_control_daemon_CP_8401_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= vector_control_daemon_CP_8401_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  vector_control_daemon_CP_8401: Block -- control-path 
    signal cp_elements: BooleanArray(2169 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= vector_control_daemon_CP_8401_start;
    vector_control_daemon_CP_8401_symbol <= cp_elements(1);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 1075 
    -- members (4) 
      -- 	$entry
      -- 	branch_block_stmt_1659/$entry
      -- 	branch_block_stmt_1659/branch_block_stmt_1659__entry__
      -- 	branch_block_stmt_1659/bb_0_bb_1
      -- 
    -- CP-element group 1 transition  place  bypass 
    -- predecessors 
    -- successors 
    -- members (3) 
      -- 	$exit
      -- 	branch_block_stmt_1659/$exit
      -- 	branch_block_stmt_1659/branch_block_stmt_1659__exit__
      -- 
    cp_elements(1) <= false; 
    -- CP-element group 2 place  bypass 
    -- predecessors 1169 
    -- successors 63 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1661__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1721__entry__
      -- 
    cp_elements(2) <= cp_elements(1169);
    -- CP-element group 3 merge  place  bypass 
    -- predecessors 95 99 
    -- successors 102 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1745__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760__entry__
      -- 
    cp_elements(3) <= OrReduce(cp_elements(95) & cp_elements(99));
    -- CP-element group 4 merge  place  bypass 
    -- predecessors 120 124 
    -- successors 127 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1774__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788__entry__
      -- 
    cp_elements(4) <= OrReduce(cp_elements(120) & cp_elements(124));
    -- CP-element group 5 merge  place  bypass 
    -- predecessors 172 178 
    -- successors 179 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1848__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1854__entry__
      -- 
    cp_elements(5) <= OrReduce(cp_elements(172) & cp_elements(178));
    -- CP-element group 6 merge  fork  transition  place  bypass 
    -- predecessors 184 190 
    -- successors 1224 1226 
    -- members (7) 
      -- 	branch_block_stmt_1659/merge_stmt_1861__exit__
      -- 	branch_block_stmt_1659/bb_7_bb_8
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$entry
      -- 
    cp_elements(6) <= OrReduce(cp_elements(184) & cp_elements(190));
    -- CP-element group 7 merge  place  bypass 
    -- predecessors 204 210 
    -- successors 211 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1898__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1904__entry__
      -- 
    cp_elements(7) <= OrReduce(cp_elements(204) & cp_elements(210));
    -- CP-element group 8 merge  place  bypass 
    -- predecessors 216 222 
    -- successors 223 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_1911__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1917__entry__
      -- 
    cp_elements(8) <= OrReduce(cp_elements(216) & cp_elements(222));
    -- CP-element group 9 branch  place  bypass 
    -- predecessors 253 
    -- successors 254 255 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_1962__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961__exit__
      -- 
    cp_elements(9) <= cp_elements(253);
    -- CP-element group 10 merge  place  bypass 
    -- predecessors 254 260 
    -- successors 261 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044__entry__
      -- 	branch_block_stmt_1659/merge_stmt_1968__exit__
      -- 
    cp_elements(10) <= OrReduce(cp_elements(254) & cp_elements(260));
    -- CP-element group 11 branch  place  bypass 
    -- predecessors 309 
    -- successors 310 311 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044__exit__
      -- 
    cp_elements(11) <= cp_elements(309);
    -- CP-element group 12 merge  place  bypass 
    -- predecessors 310 332 
    -- successors 1246 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2055__exit__
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5
      -- 
    cp_elements(12) <= OrReduce(cp_elements(310) & cp_elements(332));
    -- CP-element group 13 place  bypass 
    -- predecessors 1288 
    -- successors 333 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2057__exit__
      -- 
    cp_elements(13) <= cp_elements(1288);
    -- CP-element group 14 merge  place  bypass 
    -- predecessors 343 347 
    -- successors 1309 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2089__exit__
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8
      -- 
    cp_elements(14) <= OrReduce(cp_elements(343) & cp_elements(347));
    -- CP-element group 15 place  bypass 
    -- predecessors 1331 
    -- successors 350 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2091__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122__entry__
      -- 
    cp_elements(15) <= cp_elements(1331);
    -- CP-element group 16 branch  place  bypass 
    -- predecessors 364 
    -- successors 365 366 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_2123__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122__exit__
      -- 
    cp_elements(16) <= cp_elements(364);
    -- CP-element group 17 merge  place  bypass 
    -- predecessors 365 1350 
    -- successors 1369 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2129__exit__
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11
      -- 
    cp_elements(17) <= OrReduce(cp_elements(365) & cp_elements(1350));
    -- CP-element group 18 place  bypass 
    -- predecessors 1393 
    -- successors 372 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2140__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169__entry__
      -- 
    cp_elements(18) <= cp_elements(1393);
    -- CP-element group 19 branch  place  bypass 
    -- predecessors 390 
    -- successors 391 392 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_2170__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169__exit__
      -- 
    cp_elements(19) <= cp_elements(390);
    -- CP-element group 20 merge  fork  transition  place  bypass 
    -- predecessors 391 1399 
    -- successors 1403 1405 
    -- members (7) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13
      -- 	branch_block_stmt_1659/merge_stmt_2176__exit__
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/$entry
      -- 
    cp_elements(20) <= OrReduce(cp_elements(391) & cp_elements(1399));
    -- CP-element group 21 merge  place  bypass 
    -- predecessors 416 420 
    -- successors 1456 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20
      -- 	branch_block_stmt_1659/merge_stmt_2232__exit__
      -- 
    cp_elements(21) <= OrReduce(cp_elements(416) & cp_elements(420));
    -- CP-element group 22 place  bypass 
    -- predecessors 1478 
    -- successors 423 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2234__exit__
      -- 
    cp_elements(22) <= cp_elements(1478);
    -- CP-element group 23 branch  place  bypass 
    -- predecessors 449 
    -- successors 450 451 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_2286__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285__exit__
      -- 
    cp_elements(23) <= cp_elements(449);
    -- CP-element group 24 merge  place  bypass 
    -- predecessors 450 1497 
    -- successors 457 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2292__exit__
      -- 
    cp_elements(24) <= OrReduce(cp_elements(450) & cp_elements(1497));
    -- CP-element group 25 place  bypass 
    -- predecessors 1554 
    -- successors 475 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2325__exit__
      -- 
    cp_elements(25) <= cp_elements(1554);
    -- CP-element group 26 branch  place  bypass 
    -- predecessors 522 
    -- successors 523 524 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_2407__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406__exit__
      -- 
    cp_elements(26) <= cp_elements(522);
    -- CP-element group 27 merge  place  bypass 
    -- predecessors 523 529 
    -- successors 530 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2413__exit__
      -- 
    cp_elements(27) <= OrReduce(cp_elements(523) & cp_elements(529));
    -- CP-element group 28 branch  place  bypass 
    -- predecessors 578 
    -- successors 579 580 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489__exit__
      -- 
    cp_elements(28) <= cp_elements(578);
    -- CP-element group 29 merge  place  bypass 
    -- predecessors 579 601 
    -- successors 1566 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_2500__exit__
      -- 
    cp_elements(29) <= OrReduce(cp_elements(579) & cp_elements(601));
    -- CP-element group 30 place  bypass 
    -- predecessors 1608 
    -- successors 602 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2502__exit__
      -- 
    cp_elements(30) <= cp_elements(1608);
    -- CP-element group 31 merge  place  bypass 
    -- predecessors 612 616 
    -- successors 1629 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_2534__exit__
      -- 
    cp_elements(31) <= OrReduce(cp_elements(612) & cp_elements(616));
    -- CP-element group 32 place  bypass 
    -- predecessors 1651 
    -- successors 619 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2536__exit__
      -- 
    cp_elements(32) <= cp_elements(1651);
    -- CP-element group 33 branch  place  bypass 
    -- predecessors 633 
    -- successors 634 635 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567__exit__
      -- 	branch_block_stmt_1659/if_stmt_2568__entry__
      -- 
    cp_elements(33) <= cp_elements(633);
    -- CP-element group 34 merge  place  bypass 
    -- predecessors 634 1670 
    -- successors 1689 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_2574__exit__
      -- 
    cp_elements(34) <= OrReduce(cp_elements(634) & cp_elements(1670));
    -- CP-element group 35 place  bypass 
    -- predecessors 1713 
    -- successors 641 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2585__exit__
      -- 
    cp_elements(35) <= cp_elements(1713);
    -- CP-element group 36 branch  place  bypass 
    -- predecessors 659 
    -- successors 660 661 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614__exit__
      -- 	branch_block_stmt_1659/if_stmt_2615__entry__
      -- 
    cp_elements(36) <= cp_elements(659);
    -- CP-element group 37 merge  fork  transition  place  bypass 
    -- predecessors 660 1719 
    -- successors 1723 1725 
    -- members (7) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_2621__exit__
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/$entry
      -- 
    cp_elements(37) <= OrReduce(cp_elements(660) & cp_elements(1719));
    -- CP-element group 38 merge  place  bypass 
    -- predecessors 685 689 
    -- successors 1776 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2677__exit__
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi
      -- 
    cp_elements(38) <= OrReduce(cp_elements(685) & cp_elements(689));
    -- CP-element group 39 place  bypass 
    -- predecessors 1798 
    -- successors 692 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2679__exit__
      -- 
    cp_elements(39) <= cp_elements(1798);
    -- CP-element group 40 branch  place  bypass 
    -- predecessors 718 
    -- successors 719 720 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730__exit__
      -- 	branch_block_stmt_1659/if_stmt_2731__entry__
      -- 
    cp_elements(40) <= cp_elements(718);
    -- CP-element group 41 merge  place  bypass 
    -- predecessors 719 1817 
    -- successors 726 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2737__exit__
      -- 
    cp_elements(41) <= OrReduce(cp_elements(719) & cp_elements(1817));
    -- CP-element group 42 place  bypass 
    -- predecessors 1874 
    -- successors 744 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2770__exit__
      -- 
    cp_elements(42) <= cp_elements(1874);
    -- CP-element group 43 merge  place  bypass 
    -- predecessors 795 801 
    -- successors 802 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2878__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2872__exit__
      -- 
    cp_elements(43) <= OrReduce(cp_elements(795) & cp_elements(801));
    -- CP-element group 44 merge  fork  transition  place  bypass 
    -- predecessors 807 813 
    -- successors 1889 1891 
    -- members (7) 
      -- 	branch_block_stmt_1659/bb_43_bb_44
      -- 	branch_block_stmt_1659/merge_stmt_2885__exit__
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$entry
      -- 
    cp_elements(44) <= OrReduce(cp_elements(807) & cp_elements(813));
    -- CP-element group 45 merge  place  bypass 
    -- predecessors 827 833 
    -- successors 834 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2928__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2922__exit__
      -- 
    cp_elements(45) <= OrReduce(cp_elements(827) & cp_elements(833));
    -- CP-element group 46 merge  place  bypass 
    -- predecessors 839 845 
    -- successors 846 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2941__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2935__exit__
      -- 
    cp_elements(46) <= OrReduce(cp_elements(839) & cp_elements(845));
    -- CP-element group 47 merge  place  bypass 
    -- predecessors 851 1913 
    -- successors 858 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2948__exit__
      -- 
    cp_elements(47) <= OrReduce(cp_elements(851) & cp_elements(1913));
    -- CP-element group 48 place  bypass 
    -- predecessors 1956 
    -- successors 872 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2983__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009__entry__
      -- 
    cp_elements(48) <= cp_elements(1956);
    -- CP-element group 49 merge  place  bypass 
    -- predecessors 880 884 
    -- successors 1971 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_3016__exit__
      -- 
    cp_elements(49) <= OrReduce(cp_elements(880) & cp_elements(884));
    -- CP-element group 50 place  bypass 
    -- predecessors 1985 
    -- successors 887 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_3018__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050__entry__
      -- 
    cp_elements(50) <= cp_elements(1985);
    -- CP-element group 51 branch  place  bypass 
    -- predecessors 901 
    -- successors 902 903 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_3051__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050__exit__
      -- 
    cp_elements(51) <= cp_elements(901);
    -- CP-element group 52 merge  place  bypass 
    -- predecessors 902 2004 
    -- successors 2015 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_3057__exit__
      -- 
    cp_elements(52) <= OrReduce(cp_elements(902) & cp_elements(2004));
    -- CP-element group 53 place  bypass 
    -- predecessors 2033 
    -- successors 909 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3068__exit__
      -- 
    cp_elements(53) <= cp_elements(2033);
    -- CP-element group 54 branch  place  bypass 
    -- predecessors 925 
    -- successors 926 927 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_3100__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099__exit__
      -- 
    cp_elements(54) <= cp_elements(925);
    -- CP-element group 55 merge  place  bypass 
    -- predecessors 926 2039 
    -- successors 933 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3106__exit__
      -- 
    cp_elements(55) <= OrReduce(cp_elements(926) & cp_elements(2039));
    -- CP-element group 56 branch  place  bypass 
    -- predecessors 965 
    -- successors 966 967 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_3161__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160__exit__
      -- 
    cp_elements(56) <= cp_elements(965);
    -- CP-element group 57 merge  place  bypass 
    -- predecessors 966 970 
    -- successors 2060 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi
      -- 	branch_block_stmt_1659/merge_stmt_3167__exit__
      -- 
    cp_elements(57) <= OrReduce(cp_elements(966) & cp_elements(970));
    -- CP-element group 58 place  bypass 
    -- predecessors 2082 
    -- successors 973 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3169__exit__
      -- 
    cp_elements(58) <= cp_elements(2082);
    -- CP-element group 59 branch  place  bypass 
    -- predecessors 999 
    -- successors 1000 1001 
    -- members (2) 
      -- 	branch_block_stmt_1659/if_stmt_3221__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220__exit__
      -- 
    cp_elements(59) <= cp_elements(999);
    -- CP-element group 60 merge  place  bypass 
    -- predecessors 1000 2101 
    -- successors 1007 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3227__exit__
      -- 
    cp_elements(60) <= OrReduce(cp_elements(1000) & cp_elements(2101));
    -- CP-element group 61 place  bypass 
    -- predecessors 2158 
    -- successors 1017 
    -- members (2) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3249__exit__
      -- 
    cp_elements(61) <= cp_elements(2158);
    -- CP-element group 62 place  bypass 
    -- predecessors 1074 
    -- successors 1109 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334__exit__
      -- 
    cp_elements(62) <= cp_elements(1074);
    -- CP-element group 63 fork  transition  bypass 
    -- predecessors 2 
    -- successors 64 65 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1721/$entry
      -- 
    cp_elements(63) <= cp_elements(2);
    -- CP-element group 64 transition  output  bypass 
    -- predecessors 63 
    -- successors 66 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Sample/rr
      -- 
    cp_elements(64) <= cp_elements(63);
    rr_8696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => RPIPE_in_data_1720_inst_req_0); -- 
    -- CP-element group 65 transition  output  bypass 
    -- predecessors 63 
    -- successors 67 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Update/cr
      -- 
    cp_elements(65) <= cp_elements(63);
    cr_8701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => RPIPE_in_data_1720_inst_req_1); -- 
    -- CP-element group 66 transition  input  bypass 
    -- predecessors 64 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Sample/ra
      -- 
    ra_8697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1720_inst_ack_0, ack => cp_elements(66)); -- 
    -- CP-element group 67 transition  place  input  bypass 
    -- predecessors 65 
    -- successors 68 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1721__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1724__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1721/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1721/RPIPE_in_data_1720_Update/ca
      -- 
    ca_8702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1720_inst_ack_1, ack => cp_elements(67)); -- 
    -- CP-element group 68 fork  transition  bypass 
    -- predecessors 67 
    -- successors 69 70 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1724/$entry
      -- 
    cp_elements(68) <= cp_elements(67);
    -- CP-element group 69 transition  output  bypass 
    -- predecessors 68 
    -- successors 71 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Sample/rr
      -- 
    cp_elements(69) <= cp_elements(68);
    rr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => RPIPE_in_data_1723_inst_req_0); -- 
    -- CP-element group 70 transition  output  bypass 
    -- predecessors 68 
    -- successors 72 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Update/cr
      -- 
    cp_elements(70) <= cp_elements(68);
    cr_8718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => RPIPE_in_data_1723_inst_req_1); -- 
    -- CP-element group 71 transition  input  bypass 
    -- predecessors 69 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Sample/ra
      -- 
    ra_8714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1723_inst_ack_0, ack => cp_elements(71)); -- 
    -- CP-element group 72 transition  place  input  bypass 
    -- predecessors 70 
    -- successors 73 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1724__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1727__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1724/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1724/RPIPE_in_data_1723_Update/ca
      -- 
    ca_8719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1723_inst_ack_1, ack => cp_elements(72)); -- 
    -- CP-element group 73 fork  transition  bypass 
    -- predecessors 72 
    -- successors 74 75 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1727/$entry
      -- 
    cp_elements(73) <= cp_elements(72);
    -- CP-element group 74 transition  output  bypass 
    -- predecessors 73 
    -- successors 76 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Sample/rr
      -- 
    cp_elements(74) <= cp_elements(73);
    rr_8730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => RPIPE_in_data_1726_inst_req_0); -- 
    -- CP-element group 75 transition  output  bypass 
    -- predecessors 73 
    -- successors 77 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Update/cr
      -- 
    cp_elements(75) <= cp_elements(73);
    cr_8735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => RPIPE_in_data_1726_inst_req_1); -- 
    -- CP-element group 76 transition  input  bypass 
    -- predecessors 74 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Sample/ra
      -- 
    ra_8731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1726_inst_ack_0, ack => cp_elements(76)); -- 
    -- CP-element group 77 transition  place  input  bypass 
    -- predecessors 75 
    -- successors 78 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1727__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1730__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1727/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1727/RPIPE_in_data_1726_Update/ca
      -- 
    ca_8736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1726_inst_ack_1, ack => cp_elements(77)); -- 
    -- CP-element group 78 fork  transition  bypass 
    -- predecessors 77 
    -- successors 79 80 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1730/$entry
      -- 
    cp_elements(78) <= cp_elements(77);
    -- CP-element group 79 transition  output  bypass 
    -- predecessors 78 
    -- successors 81 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Sample/rr
      -- 
    cp_elements(79) <= cp_elements(78);
    rr_8747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => RPIPE_in_data_1729_inst_req_0); -- 
    -- CP-element group 80 transition  output  bypass 
    -- predecessors 78 
    -- successors 82 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Update/cr
      -- 
    cp_elements(80) <= cp_elements(78);
    cr_8752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => RPIPE_in_data_1729_inst_req_1); -- 
    -- CP-element group 81 transition  input  bypass 
    -- predecessors 79 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Sample/ra
      -- 
    ra_8748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1729_inst_ack_0, ack => cp_elements(81)); -- 
    -- CP-element group 82 transition  place  input  bypass 
    -- predecessors 80 
    -- successors 83 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1730__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1733__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1730/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1730/RPIPE_in_data_1729_Update/ca
      -- 
    ca_8753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1729_inst_ack_1, ack => cp_elements(82)); -- 
    -- CP-element group 83 fork  transition  bypass 
    -- predecessors 82 
    -- successors 84 85 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1733/$entry
      -- 
    cp_elements(83) <= cp_elements(82);
    -- CP-element group 84 transition  output  bypass 
    -- predecessors 83 
    -- successors 86 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Sample/rr
      -- 
    cp_elements(84) <= cp_elements(83);
    rr_8764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => RPIPE_in_data_1732_inst_req_0); -- 
    -- CP-element group 85 transition  output  bypass 
    -- predecessors 83 
    -- successors 87 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Update/cr
      -- 
    cp_elements(85) <= cp_elements(83);
    cr_8769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => RPIPE_in_data_1732_inst_req_1); -- 
    -- CP-element group 86 transition  input  bypass 
    -- predecessors 84 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Sample/ra
      -- 
    ra_8765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1732_inst_ack_0, ack => cp_elements(86)); -- 
    -- CP-element group 87 transition  place  input  bypass 
    -- predecessors 85 
    -- successors 88 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1733__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1738__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1733/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1733/RPIPE_in_data_1732_Update/ca
      -- 
    ca_8770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1732_inst_ack_1, ack => cp_elements(87)); -- 
    -- CP-element group 88 fork  transition  bypass 
    -- predecessors 87 
    -- successors 90 91 92 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/$entry
      -- 
    cp_elements(88) <= cp_elements(87);
    -- CP-element group 89 join  transition  output  bypass 
    -- predecessors 91 92 
    -- successors 93 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Sample/rr
      -- 
    cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 19) := "cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(91) & cp_elements(92);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(89), clk => clk, reset => reset); --
    end block;
    rr_8789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => SLT_f32_u1_1737_inst_req_0); -- 
    -- CP-element group 90 transition  output  bypass 
    -- predecessors 88 
    -- successors 94 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Update/cr
      -- 
    cp_elements(90) <= cp_elements(88);
    cr_8794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => SLT_f32_u1_1737_inst_req_1); -- 
    -- CP-element group 91 transition  bypass 
    -- predecessors 88 
    -- successors 89 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_speed_refx_x1_1735_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_speed_refx_x1_1735_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_speed_refx_x1_1735_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_speed_refx_x1_1735_update_completed_
      -- 
    cp_elements(91) <= cp_elements(88);
    -- CP-element group 92 transition  bypass 
    -- predecessors 88 
    -- successors 89 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_iNsTr_8_1736_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_iNsTr_8_1736_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_iNsTr_8_1736_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1738/R_iNsTr_8_1736_update_completed_
      -- 
    cp_elements(92) <= cp_elements(88);
    -- CP-element group 93 transition  input  bypass 
    -- predecessors 89 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Sample/ra
      -- 
    ra_8790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_1737_inst_ack_0, ack => cp_elements(93)); -- 
    -- CP-element group 94 branch  transition  place  input  bypass 
    -- predecessors 90 
    -- successors 95 96 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1738__exit__
      -- 	branch_block_stmt_1659/if_stmt_1739__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1738/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1738/SLT_f32_u1_1737_Update/ca
      -- 
    ca_8795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_1737_inst_ack_1, ack => cp_elements(94)); -- 
    -- CP-element group 95 transition  place  dead  bypass 
    -- predecessors 94 
    -- successors 3 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1739__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1745__entry__
      -- 	branch_block_stmt_1659/if_stmt_1739_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_1739_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1739_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_1745_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1745_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1745_dead_link/dead_transition
      -- 
    cp_elements(95) <= false;
    -- CP-element group 96 transition  output  bypass 
    -- predecessors 94 
    -- successors 97 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1739_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_1739_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1739_eval_test/branch_req
      -- 
    cp_elements(96) <= cp_elements(94);
    branch_req_8803_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => if_stmt_1739_branch_req_0); -- 
    -- CP-element group 97 branch  place  bypass 
    -- predecessors 96 
    -- successors 98 100 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_11_1740_place
      -- 
    cp_elements(97) <= cp_elements(96);
    -- CP-element group 98 transition  bypass 
    -- predecessors 97 
    -- successors 99 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1739_if_link/$entry
      -- 
    cp_elements(98) <= cp_elements(97);
    -- CP-element group 99 transition  place  input  bypass 
    -- predecessors 98 
    -- successors 3 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1739_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1739_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_1_bb_2
      -- 	branch_block_stmt_1659/merge_stmt_1745_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_1_bb_2_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_1_bb_2_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1745_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1745_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1745_PhiAck/dummy
      -- 
    if_choice_transition_8808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1739_branch_ack_1, ack => cp_elements(99)); -- 
    -- CP-element group 100 transition  bypass 
    -- predecessors 97 
    -- successors 101 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1739_else_link/$entry
      -- 
    cp_elements(100) <= cp_elements(97);
    -- CP-element group 101 transition  place  input  bypass 
    -- predecessors 100 
    -- successors 113 
    -- members (11) 
      -- 	branch_block_stmt_1659/merge_stmt_1762__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1767__entry__
      -- 	branch_block_stmt_1659/if_stmt_1739_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1739_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_1_bb_3
      -- 	branch_block_stmt_1659/merge_stmt_1762_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_1_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_1_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1762_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1762_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1762_PhiAck/dummy
      -- 
    else_choice_transition_8812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1739_branch_ack_0, ack => cp_elements(101)); -- 
    -- CP-element group 102 fork  transition  bypass 
    -- predecessors 3 
    -- successors 103 104 107 110 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/$entry
      -- 
    cp_elements(102) <= cp_elements(3);
    -- CP-element group 103 transition  output  bypass 
    -- predecessors 102 
    -- successors 106 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Update/cr
      -- 
    cp_elements(103) <= cp_elements(102);
    cr_8834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => type_cast_1749_inst_req_1); -- 
    -- CP-element group 104 transition  output  bypass 
    -- predecessors 102 
    -- successors 105 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_speed_refx_x1_1748_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_speed_refx_x1_1748_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_speed_refx_x1_1748_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_speed_refx_x1_1748_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Sample/rr
      -- 
    cp_elements(104) <= cp_elements(102);
    rr_8829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => type_cast_1749_inst_req_0); -- 
    -- CP-element group 105 transition  input  bypass 
    -- predecessors 104 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Sample/ra
      -- 
    ra_8830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_0, ack => cp_elements(105)); -- 
    -- CP-element group 106 transition  input  output  bypass 
    -- predecessors 103 
    -- successors 108 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1749_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_13_1752_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_13_1752_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_13_1752_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_13_1752_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Sample/rr
      -- 
    ca_8835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_1, ack => cp_elements(106)); -- 
    rr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ADD_f64_f64_1755_inst_req_0); -- 
    -- CP-element group 107 transition  output  bypass 
    -- predecessors 102 
    -- successors 109 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Update/cr
      -- 
    cp_elements(107) <= cp_elements(102);
    cr_8852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ADD_f64_f64_1755_inst_req_1); -- 
    -- CP-element group 108 transition  input  bypass 
    -- predecessors 106 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Sample/ra
      -- 
    ra_8848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f64_f64_1755_inst_ack_0, ack => cp_elements(108)); -- 
    -- CP-element group 109 transition  input  output  bypass 
    -- predecessors 107 
    -- successors 111 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/ADD_f64_f64_1755_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_14_1758_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_14_1758_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_14_1758_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/R_iNsTr_14_1758_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Sample/rr
      -- 
    ca_8853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f64_f64_1755_inst_ack_1, ack => cp_elements(109)); -- 
    rr_8865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => type_cast_1759_inst_req_0); -- 
    -- CP-element group 110 transition  output  bypass 
    -- predecessors 102 
    -- successors 112 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Update/cr
      -- 
    cp_elements(110) <= cp_elements(102);
    cr_8870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => type_cast_1759_inst_req_1); -- 
    -- CP-element group 111 transition  input  bypass 
    -- predecessors 109 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Sample/ra
      -- 
    ra_8866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_0, ack => cp_elements(111)); -- 
    -- CP-element group 112 fork  transition  place  input  bypass 
    -- predecessors 110 
    -- successors 1170 1176 1180 
    -- members (9) 
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760__exit__
      -- 	branch_block_stmt_1659/bb_2_bb_5
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1750_to_assign_stmt_1760/type_cast_1759_Update/ca
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$entry
      -- 
    ca_8871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_1, ack => cp_elements(112)); -- 
    -- CP-element group 113 fork  transition  bypass 
    -- predecessors 101 
    -- successors 115 116 117 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/$entry
      -- 
    cp_elements(113) <= cp_elements(101);
    -- CP-element group 114 join  transition  output  bypass 
    -- predecessors 116 117 
    -- successors 118 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Sample/rr
      -- 
    cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(116) & cp_elements(117);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(114), clk => clk, reset => reset); --
    end block;
    rr_8890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => SGT_f32_u1_1766_inst_req_0); -- 
    -- CP-element group 115 transition  output  bypass 
    -- predecessors 113 
    -- successors 119 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Update/cr
      -- 
    cp_elements(115) <= cp_elements(113);
    cr_8895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => SGT_f32_u1_1766_inst_req_1); -- 
    -- CP-element group 116 transition  bypass 
    -- predecessors 113 
    -- successors 114 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_speed_refx_x1_1764_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_speed_refx_x1_1764_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_speed_refx_x1_1764_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_speed_refx_x1_1764_update_completed_
      -- 
    cp_elements(116) <= cp_elements(113);
    -- CP-element group 117 transition  bypass 
    -- predecessors 113 
    -- successors 114 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_iNsTr_8_1765_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_iNsTr_8_1765_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_iNsTr_8_1765_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1767/R_iNsTr_8_1765_update_completed_
      -- 
    cp_elements(117) <= cp_elements(113);
    -- CP-element group 118 transition  input  bypass 
    -- predecessors 114 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Sample/ra
      -- 
    ra_8891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_1766_inst_ack_0, ack => cp_elements(118)); -- 
    -- CP-element group 119 branch  transition  place  input  bypass 
    -- predecessors 115 
    -- successors 120 121 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1767__exit__
      -- 	branch_block_stmt_1659/if_stmt_1768__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1767/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1767/SGT_f32_u1_1766_Update/ca
      -- 
    ca_8896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_1766_inst_ack_1, ack => cp_elements(119)); -- 
    -- CP-element group 120 transition  place  dead  bypass 
    -- predecessors 119 
    -- successors 4 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1768__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1774__entry__
      -- 	branch_block_stmt_1659/if_stmt_1768_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_1768_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1768_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_1774_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1774_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1774_dead_link/dead_transition
      -- 
    cp_elements(120) <= false;
    -- CP-element group 121 transition  output  bypass 
    -- predecessors 119 
    -- successors 122 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1768_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_1768_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1768_eval_test/branch_req
      -- 
    cp_elements(121) <= cp_elements(119);
    branch_req_8904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => if_stmt_1768_branch_req_0); -- 
    -- CP-element group 122 branch  place  bypass 
    -- predecessors 121 
    -- successors 123 125 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_17_1769_place
      -- 
    cp_elements(122) <= cp_elements(121);
    -- CP-element group 123 transition  bypass 
    -- predecessors 122 
    -- successors 124 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1768_if_link/$entry
      -- 
    cp_elements(123) <= cp_elements(122);
    -- CP-element group 124 transition  place  input  bypass 
    -- predecessors 123 
    -- successors 4 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1768_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1768_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_3_bb_4
      -- 	branch_block_stmt_1659/merge_stmt_1774_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_3_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1774_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1774_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1774_PhiAck/dummy
      -- 
    if_choice_transition_8909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1768_branch_ack_1, ack => cp_elements(124)); -- 
    -- CP-element group 125 transition  bypass 
    -- predecessors 122 
    -- successors 126 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1768_else_link/$entry
      -- 
    cp_elements(125) <= cp_elements(122);
    -- CP-element group 126 fork  transition  place  input  bypass 
    -- predecessors 125 
    -- successors 1185 1189 1193 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_1768_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1768_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_3_bb_5
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$entry
      -- 
    else_choice_transition_8913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1768_branch_ack_0, ack => cp_elements(126)); -- 
    -- CP-element group 127 fork  transition  bypass 
    -- predecessors 4 
    -- successors 128 129 132 135 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/$entry
      -- 
    cp_elements(127) <= cp_elements(4);
    -- CP-element group 128 transition  output  bypass 
    -- predecessors 127 
    -- successors 131 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Update/cr
      -- 
    cp_elements(128) <= cp_elements(127);
    cr_8935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => type_cast_1777_inst_req_1); -- 
    -- CP-element group 129 transition  output  bypass 
    -- predecessors 127 
    -- successors 130 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_speed_refx_x1_1776_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_speed_refx_x1_1776_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_speed_refx_x1_1776_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_speed_refx_x1_1776_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Sample/rr
      -- 
    cp_elements(129) <= cp_elements(127);
    rr_8930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => type_cast_1777_inst_req_0); -- 
    -- CP-element group 130 transition  input  bypass 
    -- predecessors 129 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Sample/ra
      -- 
    ra_8931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_0, ack => cp_elements(130)); -- 
    -- CP-element group 131 transition  input  output  bypass 
    -- predecessors 128 
    -- successors 133 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1777_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_28_1780_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_28_1780_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_28_1780_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_28_1780_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Sample/rr
      -- 
    ca_8936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_1, ack => cp_elements(131)); -- 
    rr_8948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ADD_f64_f64_1783_inst_req_0); -- 
    -- CP-element group 132 transition  output  bypass 
    -- predecessors 127 
    -- successors 134 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Update/cr
      -- 
    cp_elements(132) <= cp_elements(127);
    cr_8953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ADD_f64_f64_1783_inst_req_1); -- 
    -- CP-element group 133 transition  input  bypass 
    -- predecessors 131 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Sample/ra
      -- 
    ra_8949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f64_f64_1783_inst_ack_0, ack => cp_elements(133)); -- 
    -- CP-element group 134 transition  input  output  bypass 
    -- predecessors 132 
    -- successors 136 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/ADD_f64_f64_1783_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_29_1786_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_29_1786_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_29_1786_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/R_iNsTr_29_1786_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Sample/rr
      -- 
    ca_8954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f64_f64_1783_inst_ack_1, ack => cp_elements(134)); -- 
    rr_8966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => type_cast_1787_inst_req_0); -- 
    -- CP-element group 135 transition  output  bypass 
    -- predecessors 127 
    -- successors 137 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Update/cr
      -- 
    cp_elements(135) <= cp_elements(127);
    cr_8971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => type_cast_1787_inst_req_1); -- 
    -- CP-element group 136 transition  input  bypass 
    -- predecessors 134 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Sample/ra
      -- 
    ra_8967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1787_inst_ack_0, ack => cp_elements(136)); -- 
    -- CP-element group 137 fork  transition  place  input  bypass 
    -- predecessors 135 
    -- successors 1200 1204 1210 
    -- members (9) 
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788__exit__
      -- 	branch_block_stmt_1659/bb_4_bb_5
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1778_to_assign_stmt_1788/type_cast_1787_Update/ca
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$entry
      -- 
    ca_8972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1787_inst_ack_1, ack => cp_elements(137)); -- 
    -- CP-element group 138 fork  transition  bypass 
    -- predecessors 1217 
    -- successors 139 140 144 145 149 150 154 155 158 162 163 166 169 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/$entry
      -- 
    cp_elements(138) <= cp_elements(1217);
    -- CP-element group 139 transition  output  bypass 
    -- predecessors 138 
    -- successors 142 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Update/cr
      -- 
    cp_elements(139) <= cp_elements(138);
    cr_8992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => MUL_f32_f32_1804_inst_req_1); -- 
    -- CP-element group 140 transition  output  bypass 
    -- predecessors 138 
    -- successors 141 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_6_1801_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_6_1801_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_6_1801_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_6_1801_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Sample/rr
      -- 
    cp_elements(140) <= cp_elements(138);
    rr_8987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => MUL_f32_f32_1804_inst_req_0); -- 
    -- CP-element group 141 transition  input  bypass 
    -- predecessors 140 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Sample/ra
      -- 
    ra_8988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1804_inst_ack_0, ack => cp_elements(141)); -- 
    -- CP-element group 142 transition  input  bypass 
    -- predecessors 139 
    -- successors 143 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1804_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_19_1807_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_19_1807_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_19_1807_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_19_1807_update_completed_
      -- 
    ca_8993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1804_inst_ack_1, ack => cp_elements(142)); -- 
    -- CP-element group 143 join  transition  output  bypass 
    -- predecessors 142 145 
    -- successors 146 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Sample/rr
      -- 
    cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(142) & cp_elements(145);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(143), clk => clk, reset => reset); --
    end block;
    rr_9009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => ADD_f32_f32_1809_inst_req_0); -- 
    -- CP-element group 144 transition  output  bypass 
    -- predecessors 138 
    -- successors 147 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Update/cr
      -- 
    cp_elements(144) <= cp_elements(138);
    cr_9014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ADD_f32_f32_1809_inst_req_1); -- 
    -- CP-element group 145 transition  bypass 
    -- predecessors 138 
    -- successors 143 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_spd_lpf_prevx_x0_1808_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_spd_lpf_prevx_x0_1808_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_spd_lpf_prevx_x0_1808_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_spd_lpf_prevx_x0_1808_update_completed_
      -- 
    cp_elements(145) <= cp_elements(138);
    -- CP-element group 146 transition  input  bypass 
    -- predecessors 143 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Sample/ra
      -- 
    ra_9010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1809_inst_ack_0, ack => cp_elements(146)); -- 
    -- CP-element group 147 transition  input  bypass 
    -- predecessors 144 
    -- successors 148 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1809_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_20_1813_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_20_1813_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_20_1813_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_20_1813_update_completed_
      -- 
    ca_9015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1809_inst_ack_1, ack => cp_elements(147)); -- 
    -- CP-element group 148 join  transition  output  bypass 
    -- predecessors 147 150 
    -- successors 151 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Sample/rr
      -- 
    cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(147) & cp_elements(150);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(148), clk => clk, reset => reset); --
    end block;
    rr_9031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => SUB_f32_f32_1814_inst_req_0); -- 
    -- CP-element group 149 transition  output  bypass 
    -- predecessors 138 
    -- successors 152 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Update/cr
      -- 
    cp_elements(149) <= cp_elements(138);
    cr_9036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => SUB_f32_f32_1814_inst_req_1); -- 
    -- CP-element group 150 transition  bypass 
    -- predecessors 138 
    -- successors 148 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_refx_x0_1812_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_refx_x0_1812_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_refx_x0_1812_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_refx_x0_1812_update_completed_
      -- 
    cp_elements(150) <= cp_elements(138);
    -- CP-element group 151 transition  input  bypass 
    -- predecessors 148 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Sample/ra
      -- 
    ra_9032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_1814_inst_ack_0, ack => cp_elements(151)); -- 
    -- CP-element group 152 transition  input  bypass 
    -- predecessors 149 
    -- successors 153 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SUB_f32_f32_1814_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_21_1817_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_21_1817_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_21_1817_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_21_1817_update_completed_
      -- 
    ca_9037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_1814_inst_ack_1, ack => cp_elements(152)); -- 
    -- CP-element group 153 join  transition  output  bypass 
    -- predecessors 152 155 
    -- successors 156 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Sample/rr
      -- 
    cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(152) & cp_elements(155);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(153), clk => clk, reset => reset); --
    end block;
    rr_9053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ADD_f32_f32_1819_inst_req_0); -- 
    -- CP-element group 154 transition  output  bypass 
    -- predecessors 138 
    -- successors 157 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Update/cr
      -- 
    cp_elements(154) <= cp_elements(138);
    cr_9058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => ADD_f32_f32_1819_inst_req_1); -- 
    -- CP-element group 155 transition  bypass 
    -- predecessors 138 
    -- successors 153 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_err_prevx_x0_1818_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_err_prevx_x0_1818_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_err_prevx_x0_1818_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_speed_err_prevx_x0_1818_update_completed_
      -- 
    cp_elements(155) <= cp_elements(138);
    -- CP-element group 156 transition  input  bypass 
    -- predecessors 153 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Sample/ra
      -- 
    ra_9054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1819_inst_ack_0, ack => cp_elements(156)); -- 
    -- CP-element group 157 transition  input  output  bypass 
    -- predecessors 154 
    -- successors 159 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1819_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_22_1822_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_22_1822_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_22_1822_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_22_1822_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Sample/rr
      -- 
    ca_9059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1819_inst_ack_1, ack => cp_elements(157)); -- 
    rr_9071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => MUL_f32_f32_1825_inst_req_0); -- 
    -- CP-element group 158 transition  output  bypass 
    -- predecessors 138 
    -- successors 160 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Update/cr
      -- 
    cp_elements(158) <= cp_elements(138);
    cr_9076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => MUL_f32_f32_1825_inst_req_1); -- 
    -- CP-element group 159 transition  input  bypass 
    -- predecessors 157 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Sample/ra
      -- 
    ra_9072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1825_inst_ack_0, ack => cp_elements(159)); -- 
    -- CP-element group 160 transition  input  bypass 
    -- predecessors 158 
    -- successors 161 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/MUL_f32_f32_1825_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_23_1828_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_23_1828_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_23_1828_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_23_1828_update_completed_
      -- 
    ca_9077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1825_inst_ack_1, ack => cp_elements(160)); -- 
    -- CP-element group 161 join  transition  output  bypass 
    -- predecessors 160 163 
    -- successors 164 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Sample/rr
      -- 
    cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(160) & cp_elements(163);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(161), clk => clk, reset => reset); --
    end block;
    rr_9093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => ADD_f32_f32_1830_inst_req_0); -- 
    -- CP-element group 162 transition  output  bypass 
    -- predecessors 138 
    -- successors 165 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Update/cr
      -- 
    cp_elements(162) <= cp_elements(138);
    cr_9098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => ADD_f32_f32_1830_inst_req_1); -- 
    -- CP-element group 163 transition  bypass 
    -- predecessors 138 
    -- successors 161 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_int_speed_err_prevx_x0_1829_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_int_speed_err_prevx_x0_1829_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_int_speed_err_prevx_x0_1829_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_int_speed_err_prevx_x0_1829_update_completed_
      -- 
    cp_elements(163) <= cp_elements(138);
    -- CP-element group 164 transition  input  bypass 
    -- predecessors 161 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Sample/ra
      -- 
    ra_9094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1830_inst_ack_0, ack => cp_elements(164)); -- 
    -- CP-element group 165 transition  input  output  bypass 
    -- predecessors 162 
    -- successors 167 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/ADD_f32_f32_1830_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_24_1833_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_24_1833_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_24_1833_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_24_1833_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Sample/rr
      -- 
    ca_9099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1830_inst_ack_1, ack => cp_elements(165)); -- 
    rr_9111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => type_cast_1834_inst_req_0); -- 
    -- CP-element group 166 transition  output  bypass 
    -- predecessors 138 
    -- successors 168 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Update/cr
      -- 
    cp_elements(166) <= cp_elements(138);
    cr_9116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => type_cast_1834_inst_req_1); -- 
    -- CP-element group 167 transition  input  bypass 
    -- predecessors 165 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Sample/ra
      -- 
    ra_9112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1834_inst_ack_0, ack => cp_elements(167)); -- 
    -- CP-element group 168 transition  input  output  bypass 
    -- predecessors 166 
    -- successors 170 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/type_cast_1834_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_25_1837_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_25_1837_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_25_1837_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/R_iNsTr_25_1837_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Sample/rr
      -- 
    ca_9117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1834_inst_ack_1, ack => cp_elements(168)); -- 
    rr_9129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => SLT_f64_u1_1840_inst_req_0); -- 
    -- CP-element group 169 transition  output  bypass 
    -- predecessors 138 
    -- successors 171 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Update/cr
      -- 
    cp_elements(169) <= cp_elements(138);
    cr_9134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => SLT_f64_u1_1840_inst_req_1); -- 
    -- CP-element group 170 transition  input  bypass 
    -- predecessors 168 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Sample/ra
      -- 
    ra_9130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_1840_inst_ack_0, ack => cp_elements(170)); -- 
    -- CP-element group 171 branch  transition  place  input  bypass 
    -- predecessors 169 
    -- successors 172 173 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841__exit__
      -- 	branch_block_stmt_1659/if_stmt_1842__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841/SLT_f64_u1_1840_Update/ca
      -- 
    ca_9135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_1840_inst_ack_1, ack => cp_elements(171)); -- 
    -- CP-element group 172 transition  place  dead  bypass 
    -- predecessors 171 
    -- successors 5 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1842__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1848__entry__
      -- 	branch_block_stmt_1659/if_stmt_1842_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_1842_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1842_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_1848_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1848_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1848_dead_link/dead_transition
      -- 
    cp_elements(172) <= false;
    -- CP-element group 173 transition  output  bypass 
    -- predecessors 171 
    -- successors 174 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1842_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_1842_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1842_eval_test/branch_req
      -- 
    cp_elements(173) <= cp_elements(171);
    branch_req_9143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => if_stmt_1842_branch_req_0); -- 
    -- CP-element group 174 branch  place  bypass 
    -- predecessors 173 
    -- successors 175 177 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_26_1843_place
      -- 
    cp_elements(174) <= cp_elements(173);
    -- CP-element group 175 transition  bypass 
    -- predecessors 174 
    -- successors 176 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1842_if_link/$entry
      -- 
    cp_elements(175) <= cp_elements(174);
    -- CP-element group 176 fork  transition  place  input  bypass 
    -- predecessors 175 
    -- successors 1218 1219 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1842_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1842_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_5_bb_8
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$entry
      -- 
    if_choice_transition_9148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1842_branch_ack_1, ack => cp_elements(176)); -- 
    -- CP-element group 177 transition  bypass 
    -- predecessors 174 
    -- successors 178 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1842_else_link/$entry
      -- 
    cp_elements(177) <= cp_elements(174);
    -- CP-element group 178 transition  place  input  bypass 
    -- predecessors 177 
    -- successors 5 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1842_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1842_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_5_bb_6
      -- 	branch_block_stmt_1659/merge_stmt_1848_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_5_bb_6_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_6_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1848_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1848_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1848_PhiAck/dummy
      -- 
    else_choice_transition_9152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1842_branch_ack_0, ack => cp_elements(178)); -- 
    -- CP-element group 179 fork  transition  bypass 
    -- predecessors 5 
    -- successors 180 181 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1854/$entry
      -- 
    cp_elements(179) <= cp_elements(5);
    -- CP-element group 180 transition  output  bypass 
    -- predecessors 179 
    -- successors 183 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Update/cr
      -- 
    cp_elements(180) <= cp_elements(179);
    cr_9174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => SGT_f64_u1_1853_inst_req_1); -- 
    -- CP-element group 181 transition  output  bypass 
    -- predecessors 179 
    -- successors 182 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1854/R_iNsTr_25_1850_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1854/R_iNsTr_25_1850_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1854/R_iNsTr_25_1850_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1854/R_iNsTr_25_1850_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Sample/rr
      -- 
    cp_elements(181) <= cp_elements(179);
    rr_9169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => SGT_f64_u1_1853_inst_req_0); -- 
    -- CP-element group 182 transition  input  bypass 
    -- predecessors 181 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Sample/ra
      -- 
    ra_9170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_1853_inst_ack_0, ack => cp_elements(182)); -- 
    -- CP-element group 183 branch  transition  place  input  bypass 
    -- predecessors 180 
    -- successors 184 185 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1854__exit__
      -- 	branch_block_stmt_1659/if_stmt_1855__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1854/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1854/SGT_f64_u1_1853_Update/ca
      -- 
    ca_9175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_1853_inst_ack_1, ack => cp_elements(183)); -- 
    -- CP-element group 184 transition  place  dead  bypass 
    -- predecessors 183 
    -- successors 6 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1855__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1861__entry__
      -- 	branch_block_stmt_1659/if_stmt_1855_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_1855_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1855_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_1861_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1861_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1861_dead_link/dead_transition
      -- 
    cp_elements(184) <= false;
    -- CP-element group 185 transition  output  bypass 
    -- predecessors 183 
    -- successors 186 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1855_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_1855_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1855_eval_test/branch_req
      -- 
    cp_elements(185) <= cp_elements(183);
    branch_req_9183_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => if_stmt_1855_branch_req_0); -- 
    -- CP-element group 186 branch  place  bypass 
    -- predecessors 185 
    -- successors 187 189 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_36_1856_place
      -- 
    cp_elements(186) <= cp_elements(185);
    -- CP-element group 187 transition  bypass 
    -- predecessors 186 
    -- successors 188 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1855_if_link/$entry
      -- 
    cp_elements(187) <= cp_elements(186);
    -- CP-element group 188 fork  transition  place  input  bypass 
    -- predecessors 187 
    -- successors 1221 1222 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1855_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1855_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_6_bb_8
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$entry
      -- 
    if_choice_transition_9188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1855_branch_ack_1, ack => cp_elements(188)); -- 
    -- CP-element group 189 transition  bypass 
    -- predecessors 186 
    -- successors 190 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1855_else_link/$entry
      -- 
    cp_elements(189) <= cp_elements(186);
    -- CP-element group 190 transition  place  input  bypass 
    -- predecessors 189 
    -- successors 6 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1855_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1855_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_6_bb_7
      -- 	branch_block_stmt_1659/merge_stmt_1861_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_6_bb_7_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_7_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1861_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1861_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1861_PhiAck/dummy
      -- 
    else_choice_transition_9192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1855_branch_ack_0, ack => cp_elements(190)); -- 
    -- CP-element group 191 fork  transition  bypass 
    -- predecessors 1231 
    -- successors 192 193 197 198 201 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/$entry
      -- 
    cp_elements(191) <= cp_elements(1231);
    -- CP-element group 192 transition  output  bypass 
    -- predecessors 191 
    -- successors 195 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Update/cr
      -- 
    cp_elements(192) <= cp_elements(191);
    cr_9214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => MUL_f32_f32_1879_inst_req_1); -- 
    -- CP-element group 193 transition  output  bypass 
    -- predecessors 191 
    -- successors 194 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_21_1876_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_21_1876_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_21_1876_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_21_1876_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Sample/rr
      -- 
    cp_elements(193) <= cp_elements(191);
    rr_9209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => MUL_f32_f32_1879_inst_req_0); -- 
    -- CP-element group 194 transition  input  bypass 
    -- predecessors 193 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Sample/ra
      -- 
    ra_9210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1879_inst_ack_0, ack => cp_elements(194)); -- 
    -- CP-element group 195 transition  input  bypass 
    -- predecessors 192 
    -- successors 196 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/MUL_f32_f32_1879_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_32_1883_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_32_1883_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_32_1883_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_32_1883_update_completed_
      -- 
    ca_9215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1879_inst_ack_1, ack => cp_elements(195)); -- 
    -- CP-element group 196 join  transition  output  bypass 
    -- predecessors 195 198 
    -- successors 199 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_sample_start_
      -- 
    cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(195) & cp_elements(198);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(196), clk => clk, reset => reset); --
    end block;
    rr_9231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ADD_f32_f32_1884_inst_req_0); -- 
    -- CP-element group 197 transition  output  bypass 
    -- predecessors 191 
    -- successors 200 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_update_start_
      -- 
    cp_elements(197) <= cp_elements(191);
    cr_9236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => ADD_f32_f32_1884_inst_req_1); -- 
    -- CP-element group 198 transition  bypass 
    -- predecessors 191 
    -- successors 196 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_int_speed_errx_x0_1882_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_int_speed_errx_x0_1882_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_int_speed_errx_x0_1882_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_int_speed_errx_x0_1882_update_completed_
      -- 
    cp_elements(198) <= cp_elements(191);
    -- CP-element group 199 transition  input  bypass 
    -- predecessors 196 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_sample_completed_
      -- 
    ra_9232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1884_inst_ack_0, ack => cp_elements(199)); -- 
    -- CP-element group 200 transition  input  output  bypass 
    -- predecessors 197 
    -- successors 202 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_33_1887_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_33_1887_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_33_1887_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/R_iNsTr_33_1887_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/ADD_f32_f32_1884_update_completed_
      -- 
    ca_9237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1884_inst_ack_1, ack => cp_elements(200)); -- 
    rr_9249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => SLT_f32_u1_1890_inst_req_0); -- 
    -- CP-element group 201 transition  output  bypass 
    -- predecessors 191 
    -- successors 203 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Update/$entry
      -- 
    cp_elements(201) <= cp_elements(191);
    cr_9254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => SLT_f32_u1_1890_inst_req_1); -- 
    -- CP-element group 202 transition  input  bypass 
    -- predecessors 200 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Sample/$exit
      -- 
    ra_9250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_1890_inst_ack_0, ack => cp_elements(202)); -- 
    -- CP-element group 203 branch  transition  place  input  bypass 
    -- predecessors 201 
    -- successors 204 205 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891__exit__
      -- 	branch_block_stmt_1659/if_stmt_1892__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/SLT_f32_u1_1890_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891/$exit
      -- 
    ca_9255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_1890_inst_ack_1, ack => cp_elements(203)); -- 
    -- CP-element group 204 transition  place  dead  bypass 
    -- predecessors 203 
    -- successors 7 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1892__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1898__entry__
      -- 	branch_block_stmt_1659/if_stmt_1892_dead_link/dead_transition
      -- 	branch_block_stmt_1659/if_stmt_1892_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1892_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1898_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1898_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1898_dead_link/dead_transition
      -- 
    cp_elements(204) <= false;
    -- CP-element group 205 transition  output  bypass 
    -- predecessors 203 
    -- successors 206 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1892_eval_test/branch_req
      -- 	branch_block_stmt_1659/if_stmt_1892_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1892_eval_test/$entry
      -- 
    cp_elements(205) <= cp_elements(203);
    branch_req_9263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => if_stmt_1892_branch_req_0); -- 
    -- CP-element group 206 branch  place  bypass 
    -- predecessors 205 
    -- successors 207 209 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_34_1893_place
      -- 
    cp_elements(206) <= cp_elements(205);
    -- CP-element group 207 transition  bypass 
    -- predecessors 206 
    -- successors 208 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1892_if_link/$entry
      -- 
    cp_elements(207) <= cp_elements(206);
    -- CP-element group 208 fork  transition  place  input  bypass 
    -- predecessors 207 
    -- successors 1237 1238 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1892_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/if_stmt_1892_if_link/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$entry
      -- 
    if_choice_transition_9268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1892_branch_ack_1, ack => cp_elements(208)); -- 
    -- CP-element group 209 transition  bypass 
    -- predecessors 206 
    -- successors 210 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1892_else_link/$entry
      -- 
    cp_elements(209) <= cp_elements(206);
    -- CP-element group 210 transition  place  input  bypass 
    -- predecessors 209 
    -- successors 7 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1892_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/if_stmt_1892_else_link/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_9
      -- 	branch_block_stmt_1659/bb_8_bb_9_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_9_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1898_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_1898_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1898_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1898_PhiAck/dummy
      -- 
    else_choice_transition_9272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1892_branch_ack_0, ack => cp_elements(210)); -- 
    -- CP-element group 211 fork  transition  bypass 
    -- predecessors 7 
    -- successors 212 213 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1904/$entry
      -- 
    cp_elements(211) <= cp_elements(7);
    -- CP-element group 212 transition  output  bypass 
    -- predecessors 211 
    -- successors 215 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_update_start_
      -- 
    cp_elements(212) <= cp_elements(211);
    cr_9294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => SGT_f32_u1_1903_inst_req_1); -- 
    -- CP-element group 213 transition  output  bypass 
    -- predecessors 211 
    -- successors 214 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1904/R_iNsTr_33_1900_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1904/R_iNsTr_33_1900_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1904/R_iNsTr_33_1900_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1904/R_iNsTr_33_1900_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_sample_start_
      -- 
    cp_elements(213) <= cp_elements(211);
    rr_9289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => SGT_f32_u1_1903_inst_req_0); -- 
    -- CP-element group 214 transition  input  bypass 
    -- predecessors 213 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_sample_completed_
      -- 
    ra_9290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_1903_inst_ack_0, ack => cp_elements(214)); -- 
    -- CP-element group 215 branch  transition  place  input  bypass 
    -- predecessors 212 
    -- successors 216 217 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_1904__exit__
      -- 	branch_block_stmt_1659/if_stmt_1905__entry__
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1904/SGT_f32_u1_1903_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1904/$exit
      -- 
    ca_9295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_1903_inst_ack_1, ack => cp_elements(215)); -- 
    -- CP-element group 216 transition  place  dead  bypass 
    -- predecessors 215 
    -- successors 8 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1905__exit__
      -- 	branch_block_stmt_1659/merge_stmt_1911__entry__
      -- 	branch_block_stmt_1659/if_stmt_1905_dead_link/dead_transition
      -- 	branch_block_stmt_1659/if_stmt_1905_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1905_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1911_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1911_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1911_dead_link/dead_transition
      -- 
    cp_elements(216) <= false;
    -- CP-element group 217 transition  output  bypass 
    -- predecessors 215 
    -- successors 218 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1905_eval_test/branch_req
      -- 	branch_block_stmt_1659/if_stmt_1905_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1905_eval_test/$entry
      -- 
    cp_elements(217) <= cp_elements(215);
    branch_req_9303_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => if_stmt_1905_branch_req_0); -- 
    -- CP-element group 218 branch  place  bypass 
    -- predecessors 217 
    -- successors 219 221 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_43_1906_place
      -- 
    cp_elements(218) <= cp_elements(217);
    -- CP-element group 219 transition  bypass 
    -- predecessors 218 
    -- successors 220 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1905_if_link/$entry
      -- 
    cp_elements(219) <= cp_elements(218);
    -- CP-element group 220 fork  transition  place  input  bypass 
    -- predecessors 219 
    -- successors 1240 1241 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_1905_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1905_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_9_bb_11
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$entry
      -- 
    if_choice_transition_9308_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1905_branch_ack_1, ack => cp_elements(220)); -- 
    -- CP-element group 221 transition  bypass 
    -- predecessors 218 
    -- successors 222 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1905_else_link/$entry
      -- 
    cp_elements(221) <= cp_elements(218);
    -- CP-element group 222 transition  place  input  bypass 
    -- predecessors 221 
    -- successors 8 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_1905_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1905_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_9_bb_10
      -- 	branch_block_stmt_1659/bb_9_bb_10_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_10_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1911_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_1911_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1911_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1911_PhiAck/dummy
      -- 
    else_choice_transition_9312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1905_branch_ack_0, ack => cp_elements(222)); -- 
    -- CP-element group 223 fork  transition  bypass 
    -- predecessors 8 
    -- successors 224 225 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1917/$entry
      -- 
    cp_elements(223) <= cp_elements(8);
    -- CP-element group 224 transition  output  bypass 
    -- predecessors 223 
    -- successors 227 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Update/$entry
      -- 
    cp_elements(224) <= cp_elements(223);
    cr_9334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => MUL_f32_f32_1916_inst_req_1); -- 
    -- CP-element group 225 transition  output  bypass 
    -- predecessors 223 
    -- successors 226 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1917/R_iNsTr_33_1913_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1917/R_iNsTr_33_1913_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1917/R_iNsTr_33_1913_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1917/R_iNsTr_33_1913_sample_completed_
      -- 
    cp_elements(225) <= cp_elements(223);
    rr_9329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => MUL_f32_f32_1916_inst_req_0); -- 
    -- CP-element group 226 transition  input  bypass 
    -- predecessors 225 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Sample/$exit
      -- 
    ra_9330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1916_inst_ack_0, ack => cp_elements(226)); -- 
    -- CP-element group 227 fork  transition  place  input  bypass 
    -- predecessors 224 
    -- successors 1232 1234 
    -- members (11) 
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1917/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1917__exit__
      -- 	branch_block_stmt_1659/bb_10_bb_11
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1917/MUL_f32_f32_1916_Update/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$entry
      -- 
    ca_9335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1916_inst_ack_1, ack => cp_elements(227)); -- 
    -- CP-element group 228 fork  transition  bypass 
    -- predecessors 1245 
    -- successors 229 230 234 235 238 239 242 246 249 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/$entry
      -- 
    cp_elements(228) <= cp_elements(1245);
    -- CP-element group 229 transition  output  bypass 
    -- predecessors 228 
    -- successors 232 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_update_start_
      -- 
    cp_elements(229) <= cp_elements(228);
    cr_9355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => MUL_f32_f32_1935_inst_req_1); -- 
    -- CP-element group 230 transition  output  bypass 
    -- predecessors 228 
    -- successors 231 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_2_1932_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_2_1932_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_2_1932_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_2_1932_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_sample_start_
      -- 
    cp_elements(230) <= cp_elements(228);
    rr_9350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => MUL_f32_f32_1935_inst_req_0); -- 
    -- CP-element group 231 transition  input  bypass 
    -- predecessors 230 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_sample_completed_
      -- 
    ra_9351_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1935_inst_ack_0, ack => cp_elements(231)); -- 
    -- CP-element group 232 transition  input  bypass 
    -- predecessors 229 
    -- successors 233 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_38_1938_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_38_1938_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_38_1938_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_38_1938_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1935_update_completed_
      -- 
    ca_9356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1935_inst_ack_1, ack => cp_elements(232)); -- 
    -- CP-element group 233 join  transition  output  bypass 
    -- predecessors 232 235 
    -- successors 236 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_sample_start_
      -- 
    cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(232) & cp_elements(235);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(233), clk => clk, reset => reset); --
    end block;
    rr_9372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ADD_f32_f32_1940_inst_req_0); -- 
    -- CP-element group 234 transition  output  bypass 
    -- predecessors 228 
    -- successors 237 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Update/$entry
      -- 
    cp_elements(234) <= cp_elements(228);
    cr_9377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ADD_f32_f32_1940_inst_req_1); -- 
    -- CP-element group 235 transition  bypass 
    -- predecessors 228 
    -- successors 233 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_flux_rotor_prevx_x0_1939_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_flux_rotor_prevx_x0_1939_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_flux_rotor_prevx_x0_1939_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_flux_rotor_prevx_x0_1939_update_completed_
      -- 
    cp_elements(235) <= cp_elements(228);
    -- CP-element group 236 transition  input  bypass 
    -- predecessors 233 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Sample/ra
      -- 
    ra_9373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1940_inst_ack_0, ack => cp_elements(236)); -- 
    -- CP-element group 237 transition  input  output  bypass 
    -- predecessors 234 
    -- successors 247 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_39_1953_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_39_1953_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_39_1953_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_39_1953_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/ADD_f32_f32_1940_Update/$exit
      -- 
    ca_9378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_1940_inst_ack_1, ack => cp_elements(237)); -- 
    rr_9426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => type_cast_1954_inst_req_0); -- 
    -- CP-element group 238 transition  output  bypass 
    -- predecessors 228 
    -- successors 241 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_update_start_
      -- 
    cp_elements(238) <= cp_elements(228);
    cr_9395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => MUL_f32_f32_1946_inst_req_1); -- 
    -- CP-element group 239 transition  output  bypass 
    -- predecessors 228 
    -- successors 240 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_4_1943_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_4_1943_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_4_1943_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_4_1943_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_sample_start_
      -- 
    cp_elements(239) <= cp_elements(228);
    rr_9390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => MUL_f32_f32_1946_inst_req_0); -- 
    -- CP-element group 240 transition  input  bypass 
    -- predecessors 239 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_sample_completed_
      -- 
    ra_9391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1946_inst_ack_0, ack => cp_elements(240)); -- 
    -- CP-element group 241 fork  transition  input  bypass 
    -- predecessors 238 
    -- successors 243 250 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/MUL_f32_f32_1946_update_completed_
      -- 
    ca_9396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1946_inst_ack_1, ack => cp_elements(241)); -- 
    -- CP-element group 242 transition  output  bypass 
    -- predecessors 228 
    -- successors 245 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Update/$entry
      -- 
    cp_elements(242) <= cp_elements(228);
    cr_9413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => type_cast_1950_inst_req_1); -- 
    -- CP-element group 243 transition  output  bypass 
    -- predecessors 241 
    -- successors 244 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1949_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1949_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1949_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1949_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Sample/rr
      -- 
    cp_elements(243) <= cp_elements(241);
    rr_9408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(243), ack => type_cast_1950_inst_req_0); -- 
    -- CP-element group 244 transition  input  bypass 
    -- predecessors 243 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Sample/$exit
      -- 
    ra_9409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1950_inst_ack_0, ack => cp_elements(244)); -- 
    -- CP-element group 245 transition  input  bypass 
    -- predecessors 242 
    -- successors 253 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1950_Update/$exit
      -- 
    ca_9414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1950_inst_ack_1, ack => cp_elements(245)); -- 
    -- CP-element group 246 transition  output  bypass 
    -- predecessors 228 
    -- successors 248 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Update/cr
      -- 
    cp_elements(246) <= cp_elements(228);
    cr_9431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => type_cast_1954_inst_req_1); -- 
    -- CP-element group 247 transition  input  bypass 
    -- predecessors 237 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_sample_completed_
      -- 
    ra_9427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_0, ack => cp_elements(247)); -- 
    -- CP-element group 248 transition  input  bypass 
    -- predecessors 246 
    -- successors 253 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/type_cast_1954_Update/ca
      -- 
    ca_9432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_1, ack => cp_elements(248)); -- 
    -- CP-element group 249 transition  output  bypass 
    -- predecessors 228 
    -- successors 252 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_update_start_
      -- 
    cp_elements(249) <= cp_elements(228);
    cr_9449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => EQ_f32_u1_1960_inst_req_1); -- 
    -- CP-element group 250 transition  output  bypass 
    -- predecessors 241 
    -- successors 251 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1957_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1957_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1957_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/R_iNsTr_40_1957_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_sample_start_
      -- 
    cp_elements(250) <= cp_elements(241);
    rr_9444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => EQ_f32_u1_1960_inst_req_0); -- 
    -- CP-element group 251 transition  input  bypass 
    -- predecessors 250 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_sample_completed_
      -- 
    ra_9445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_1960_inst_ack_0, ack => cp_elements(251)); -- 
    -- CP-element group 252 transition  input  bypass 
    -- predecessors 249 
    -- successors 253 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/EQ_f32_u1_1960_Update/ca
      -- 
    ca_9450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_1960_inst_ack_1, ack => cp_elements(252)); -- 
    -- CP-element group 253 join  transition  bypass 
    -- predecessors 245 248 252 
    -- successors 9 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961/$exit
      -- 
    cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(245) & cp_elements(248) & cp_elements(252);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254 transition  place  dead  bypass 
    -- predecessors 9 
    -- successors 10 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_1968__entry__
      -- 	branch_block_stmt_1659/if_stmt_1962__exit__
      -- 	branch_block_stmt_1659/if_stmt_1962_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_1962_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1962_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_1968_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1968_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1968_dead_link/dead_transition
      -- 
    cp_elements(254) <= false;
    -- CP-element group 255 transition  output  bypass 
    -- predecessors 9 
    -- successors 256 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_1962_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_1962_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_1962_eval_test/branch_req
      -- 
    cp_elements(255) <= cp_elements(9);
    branch_req_9458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => if_stmt_1962_branch_req_0); -- 
    -- CP-element group 256 branch  place  bypass 
    -- predecessors 255 
    -- successors 257 259 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_41_1963_place
      -- 
    cp_elements(256) <= cp_elements(255);
    -- CP-element group 257 transition  bypass 
    -- predecessors 256 
    -- successors 258 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1962_if_link/$entry
      -- 
    cp_elements(257) <= cp_elements(256);
    -- CP-element group 258 fork  transition  place  input  bypass 
    -- predecessors 257 
    -- successors 1555 1556 
    -- members (8) 
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit
      -- 	branch_block_stmt_1659/if_stmt_1962_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1962_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/$entry
      -- 
    if_choice_transition_9463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1962_branch_ack_1, ack => cp_elements(258)); -- 
    -- CP-element group 259 transition  bypass 
    -- predecessors 256 
    -- successors 260 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_1962_else_link/$entry
      -- 
    cp_elements(259) <= cp_elements(256);
    -- CP-element group 260 transition  place  input  bypass 
    -- predecessors 259 
    -- successors 10 
    -- members (9) 
      -- 	branch_block_stmt_1659/bb_11_bb_12
      -- 	branch_block_stmt_1659/if_stmt_1962_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_1962_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_11_bb_12_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_11_bb_12_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1968_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_1968_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_1968_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1968_PhiAck/dummy
      -- 
    else_choice_transition_9467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1962_branch_ack_0, ack => cp_elements(260)); -- 
    -- CP-element group 261 fork  transition  bypass 
    -- predecessors 10 
    -- successors 262 263 266 269 270 273 276 277 280 283 286 287 290 293 297 298 299 302 306 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/$entry
      -- 
    cp_elements(261) <= cp_elements(10);
    -- CP-element group 262 transition  output  bypass 
    -- predecessors 261 
    -- successors 265 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Update/$entry
      -- 
    cp_elements(262) <= cp_elements(261);
    cr_9489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(262), ack => LSHR_u32_u32_1973_inst_req_1); -- 
    -- CP-element group 263 transition  output  bypass 
    -- predecessors 261 
    -- successors 264 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1970_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1970_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1970_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1970_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_sample_start_
      -- 
    cp_elements(263) <= cp_elements(261);
    rr_9484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => LSHR_u32_u32_1973_inst_req_0); -- 
    -- CP-element group 264 transition  input  bypass 
    -- predecessors 263 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Sample/$exit
      -- 
    ra_9485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_1973_inst_ack_0, ack => cp_elements(264)); -- 
    -- CP-element group 265 transition  input  output  bypass 
    -- predecessors 262 
    -- successors 267 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_52_1976_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_52_1976_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_52_1976_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_52_1976_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1973_Update/$exit
      -- 
    ca_9490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_1973_inst_ack_1, ack => cp_elements(265)); -- 
    rr_9502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => AND_u32_u32_1979_inst_req_0); -- 
    -- CP-element group 266 transition  output  bypass 
    -- predecessors 261 
    -- successors 268 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_update_start_
      -- 
    cp_elements(266) <= cp_elements(261);
    cr_9507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => AND_u32_u32_1979_inst_req_1); -- 
    -- CP-element group 267 transition  input  bypass 
    -- predecessors 265 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_sample_completed_
      -- 
    ra_9503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_1979_inst_ack_0, ack => cp_elements(267)); -- 
    -- CP-element group 268 transition  input  bypass 
    -- predecessors 266 
    -- successors 305 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1979_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_53_2041_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_53_2041_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_53_2041_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_53_2041_update_completed_
      -- 
    ca_9508_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_1979_inst_ack_1, ack => cp_elements(268)); -- 
    -- CP-element group 269 transition  output  bypass 
    -- predecessors 261 
    -- successors 272 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Update/cr
      -- 
    cp_elements(269) <= cp_elements(261);
    cr_9525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => LSHR_u32_u32_1985_inst_req_1); -- 
    -- CP-element group 270 transition  output  bypass 
    -- predecessors 261 
    -- successors 271 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_1982_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_1982_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_1982_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_1982_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Sample/rr
      -- 
    cp_elements(270) <= cp_elements(261);
    rr_9520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => LSHR_u32_u32_1985_inst_req_0); -- 
    -- CP-element group 271 transition  input  bypass 
    -- predecessors 270 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Sample/ra
      -- 
    ra_9521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_1985_inst_ack_0, ack => cp_elements(271)); -- 
    -- CP-element group 272 transition  input  output  bypass 
    -- predecessors 269 
    -- successors 274 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_1985_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_54_1988_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_54_1988_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_54_1988_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_54_1988_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Sample/$entry
      -- 
    ca_9526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_1985_inst_ack_1, ack => cp_elements(272)); -- 
    rr_9538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(272), ack => AND_u32_u32_1991_inst_req_0); -- 
    -- CP-element group 273 transition  output  bypass 
    -- predecessors 261 
    -- successors 275 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Update/cr
      -- 
    cp_elements(273) <= cp_elements(261);
    cr_9543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => AND_u32_u32_1991_inst_req_1); -- 
    -- CP-element group 274 transition  input  bypass 
    -- predecessors 272 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Sample/$exit
      -- 
    ra_9539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_1991_inst_ack_0, ack => cp_elements(274)); -- 
    -- CP-element group 275 transition  input  bypass 
    -- predecessors 273 
    -- successors 305 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_1991_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_55_2042_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_55_2042_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_55_2042_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_55_2042_update_completed_
      -- 
    ca_9544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_1991_inst_ack_1, ack => cp_elements(275)); -- 
    -- CP-element group 276 transition  output  bypass 
    -- predecessors 261 
    -- successors 279 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_update_start_
      -- 
    cp_elements(276) <= cp_elements(261);
    cr_9561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => SHL_u32_u32_1997_inst_req_1); -- 
    -- CP-element group 277 transition  output  bypass 
    -- predecessors 261 
    -- successors 278 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1994_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1994_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1994_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_1994_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_sample_start_
      -- 
    cp_elements(277) <= cp_elements(261);
    rr_9556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => SHL_u32_u32_1997_inst_req_0); -- 
    -- CP-element group 278 transition  input  bypass 
    -- predecessors 277 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_sample_completed_
      -- 
    ra_9557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_1997_inst_ack_0, ack => cp_elements(278)); -- 
    -- CP-element group 279 transition  input  output  bypass 
    -- predecessors 276 
    -- successors 281 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SHL_u32_u32_1997_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_56_2000_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_56_2000_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_56_2000_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_56_2000_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Sample/rr
      -- 
    ca_9562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_1997_inst_ack_1, ack => cp_elements(279)); -- 
    rr_9574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => AND_u32_u32_2003_inst_req_0); -- 
    -- CP-element group 280 transition  output  bypass 
    -- predecessors 261 
    -- successors 282 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Update/cr
      -- 
    cp_elements(280) <= cp_elements(261);
    cr_9579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => AND_u32_u32_2003_inst_req_1); -- 
    -- CP-element group 281 transition  input  bypass 
    -- predecessors 279 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Sample/ra
      -- 
    ra_9575_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2003_inst_ack_0, ack => cp_elements(281)); -- 
    -- CP-element group 282 transition  input  output  bypass 
    -- predecessors 280 
    -- successors 284 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_57_2006_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2003_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_57_2006_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_57_2006_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_57_2006_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Sample/rr
      -- 
    ca_9580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2003_inst_ack_1, ack => cp_elements(282)); -- 
    rr_9592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => OR_u32_u32_2009_inst_req_0); -- 
    -- CP-element group 283 transition  output  bypass 
    -- predecessors 261 
    -- successors 285 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Update/cr
      -- 
    cp_elements(283) <= cp_elements(261);
    cr_9597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => OR_u32_u32_2009_inst_req_1); -- 
    -- CP-element group 284 transition  input  bypass 
    -- predecessors 282 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Sample/ra
      -- 
    ra_9593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2009_inst_ack_0, ack => cp_elements(284)); -- 
    -- CP-element group 285 transition  input  bypass 
    -- predecessors 283 
    -- successors 309 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2009_Update/ca
      -- 
    ca_9598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2009_inst_ack_1, ack => cp_elements(285)); -- 
    -- CP-element group 286 transition  output  bypass 
    -- predecessors 261 
    -- successors 289 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Update/cr
      -- 
    cp_elements(286) <= cp_elements(261);
    cr_9615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => LSHR_u32_u32_2015_inst_req_1); -- 
    -- CP-element group 287 transition  output  bypass 
    -- predecessors 261 
    -- successors 288 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2012_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2012_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2012_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2012_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Sample/rr
      -- 
    cp_elements(287) <= cp_elements(261);
    rr_9610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(287), ack => LSHR_u32_u32_2015_inst_req_0); -- 
    -- CP-element group 288 transition  input  bypass 
    -- predecessors 287 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Sample/ra
      -- 
    ra_9611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2015_inst_ack_0, ack => cp_elements(288)); -- 
    -- CP-element group 289 transition  input  output  bypass 
    -- predecessors 286 
    -- successors 291 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/LSHR_u32_u32_2015_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_59_2018_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_59_2018_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_59_2018_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_59_2018_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Sample/rr
      -- 
    ca_9616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2015_inst_ack_1, ack => cp_elements(289)); -- 
    rr_9628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => AND_u32_u32_2021_inst_req_0); -- 
    -- CP-element group 290 transition  output  bypass 
    -- predecessors 261 
    -- successors 292 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Update/cr
      -- 
    cp_elements(290) <= cp_elements(261);
    cr_9633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => AND_u32_u32_2021_inst_req_1); -- 
    -- CP-element group 291 transition  input  bypass 
    -- predecessors 289 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Sample/ra
      -- 
    ra_9629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2021_inst_ack_0, ack => cp_elements(291)); -- 
    -- CP-element group 292 transition  input  output  bypass 
    -- predecessors 290 
    -- successors 294 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2021_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_60_2024_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_60_2024_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_60_2024_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_60_2024_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Sample/rr
      -- 
    ca_9634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2021_inst_ack_1, ack => cp_elements(292)); -- 
    rr_9646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => OR_u32_u32_2027_inst_req_0); -- 
    -- CP-element group 293 transition  output  bypass 
    -- predecessors 261 
    -- successors 295 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Update/cr
      -- 
    cp_elements(293) <= cp_elements(261);
    cr_9651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => OR_u32_u32_2027_inst_req_1); -- 
    -- CP-element group 294 transition  input  bypass 
    -- predecessors 292 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Sample/ra
      -- 
    ra_9647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2027_inst_ack_0, ack => cp_elements(294)); -- 
    -- CP-element group 295 transition  input  bypass 
    -- predecessors 293 
    -- successors 309 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/OR_u32_u32_2027_Update/ca
      -- 
    ca_9652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2027_inst_ack_1, ack => cp_elements(295)); -- 
    -- CP-element group 296 join  transition  output  bypass 
    -- predecessors 298 299 
    -- successors 300 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Sample/rr
      -- 
    cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(298) & cp_elements(299);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(296), clk => clk, reset => reset); --
    end block;
    rr_9668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => XOR_u32_u32_2032_inst_req_0); -- 
    -- CP-element group 297 transition  output  bypass 
    -- predecessors 261 
    -- successors 301 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Update/cr
      -- 
    cp_elements(297) <= cp_elements(261);
    cr_9673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => XOR_u32_u32_2032_inst_req_1); -- 
    -- CP-element group 298 transition  bypass 
    -- predecessors 261 
    -- successors 296 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2030_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2030_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2030_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp6x_xix_xi2_2030_update_completed_
      -- 
    cp_elements(298) <= cp_elements(261);
    -- CP-element group 299 transition  bypass 
    -- predecessors 261 
    -- successors 296 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_2031_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_2031_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_2031_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_tmp10x_xix_xi1_2031_update_completed_
      -- 
    cp_elements(299) <= cp_elements(261);
    -- CP-element group 300 transition  input  bypass 
    -- predecessors 296 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Sample/ra
      -- 
    ra_9669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2032_inst_ack_0, ack => cp_elements(300)); -- 
    -- CP-element group 301 transition  input  output  bypass 
    -- predecessors 297 
    -- successors 303 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/XOR_u32_u32_2032_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_62_2035_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_62_2035_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_62_2035_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/R_iNsTr_62_2035_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Sample/rr
      -- 
    ca_9674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2032_inst_ack_1, ack => cp_elements(301)); -- 
    rr_9686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => AND_u32_u32_2038_inst_req_0); -- 
    -- CP-element group 302 transition  output  bypass 
    -- predecessors 261 
    -- successors 304 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Update/cr
      -- 
    cp_elements(302) <= cp_elements(261);
    cr_9691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => AND_u32_u32_2038_inst_req_1); -- 
    -- CP-element group 303 transition  input  bypass 
    -- predecessors 301 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Sample/ra
      -- 
    ra_9687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2038_inst_ack_0, ack => cp_elements(303)); -- 
    -- CP-element group 304 transition  input  bypass 
    -- predecessors 302 
    -- successors 309 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/AND_u32_u32_2038_Update/ca
      -- 
    ca_9692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2038_inst_ack_1, ack => cp_elements(304)); -- 
    -- CP-element group 305 join  transition  output  bypass 
    -- predecessors 268 275 
    -- successors 307 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Sample/rr
      -- 
    cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(268) & cp_elements(275);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(305), clk => clk, reset => reset); --
    end block;
    rr_9708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => SUB_u32_u32_2043_inst_req_0); -- 
    -- CP-element group 306 transition  output  bypass 
    -- predecessors 261 
    -- successors 308 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Update/cr
      -- 
    cp_elements(306) <= cp_elements(261);
    cr_9713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => SUB_u32_u32_2043_inst_req_1); -- 
    -- CP-element group 307 transition  input  bypass 
    -- predecessors 305 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Sample/ra
      -- 
    ra_9709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2043_inst_ack_0, ack => cp_elements(307)); -- 
    -- CP-element group 308 transition  input  bypass 
    -- predecessors 306 
    -- successors 309 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/SUB_u32_u32_2043_Update/ca
      -- 
    ca_9714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2043_inst_ack_1, ack => cp_elements(308)); -- 
    -- CP-element group 309 join  transition  bypass 
    -- predecessors 285 295 304 308 
    -- successors 11 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_1974_to_assign_stmt_2044/$exit
      -- 
    cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_309"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= cp_elements(285) & cp_elements(295) & cp_elements(304) & cp_elements(308);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310 transition  place  dead  bypass 
    -- predecessors 11 
    -- successors 12 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2055__entry__
      -- 	branch_block_stmt_1659/switch_stmt_2045__exit__
      -- 	branch_block_stmt_1659/switch_stmt_2045_dead_link/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045_dead_link/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2055_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2055_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2055_dead_link/dead_transition
      -- 
    cp_elements(310) <= false;
    -- CP-element group 311 place  bypass 
    -- predecessors 11 
    -- successors 312 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check_place__
      -- 
    cp_elements(311) <= cp_elements(11);
    -- CP-element group 312 fork  transition  bypass 
    -- predecessors 311 
    -- successors 313 319 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/$entry
      -- 
    cp_elements(312) <= cp_elements(311);
    -- CP-element group 313 fork  transition  bypass 
    -- predecessors 312 
    -- successors 314 316 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/$entry
      -- 
    cp_elements(313) <= cp_elements(312);
    -- CP-element group 314 transition  output  bypass 
    -- predecessors 313 
    -- successors 315 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Sample/rr
      -- 
    cp_elements(314) <= cp_elements(313);
    rr_9732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(314), ack => switch_stmt_2045_select_expr_0_req_0); -- 
    -- CP-element group 315 transition  input  bypass 
    -- predecessors 314 
    -- successors 318 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Sample/ra
      -- 
    ra_9733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_select_expr_0_ack_0, ack => cp_elements(315)); -- 
    -- CP-element group 316 transition  output  bypass 
    -- predecessors 313 
    -- successors 317 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Update/cr
      -- 
    cp_elements(316) <= cp_elements(313);
    cr_9737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => switch_stmt_2045_select_expr_0_req_1); -- 
    -- CP-element group 317 transition  input  bypass 
    -- predecessors 316 
    -- successors 318 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/Update/ca
      -- 
    ca_9738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_select_expr_0_ack_1, ack => cp_elements(317)); -- 
    -- CP-element group 318 join  transition  output  bypass 
    -- predecessors 315 317 
    -- successors 325 
    -- members (3) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_0/cmp
      -- 
    cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(315) & cp_elements(317);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(318), clk => clk, reset => reset); --
    end block;
    cmp_9739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => switch_stmt_2045_branch_0_req_0); -- 
    -- CP-element group 319 fork  transition  bypass 
    -- predecessors 312 
    -- successors 320 322 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/$entry
      -- 
    cp_elements(319) <= cp_elements(312);
    -- CP-element group 320 transition  output  bypass 
    -- predecessors 319 
    -- successors 321 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Sample/rr
      -- 
    cp_elements(320) <= cp_elements(319);
    rr_9749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(320), ack => switch_stmt_2045_select_expr_1_req_0); -- 
    -- CP-element group 321 transition  input  bypass 
    -- predecessors 320 
    -- successors 324 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Sample/ra
      -- 
    ra_9750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_select_expr_1_ack_0, ack => cp_elements(321)); -- 
    -- CP-element group 322 transition  output  bypass 
    -- predecessors 319 
    -- successors 323 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Update/cr
      -- 
    cp_elements(322) <= cp_elements(319);
    cr_9754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => switch_stmt_2045_select_expr_1_req_1); -- 
    -- CP-element group 323 transition  input  bypass 
    -- predecessors 322 
    -- successors 324 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/Update/ca
      -- 
    ca_9755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_select_expr_1_ack_1, ack => cp_elements(323)); -- 
    -- CP-element group 324 join  transition  output  bypass 
    -- predecessors 321 323 
    -- successors 325 
    -- members (3) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/condition_1/cmp
      -- 
    cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(321) & cp_elements(323);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(324), clk => clk, reset => reset); --
    end block;
    cmp_9756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(324), ack => switch_stmt_2045_branch_1_req_0); -- 
    -- CP-element group 325 join  transition  output  bypass 
    -- predecessors 318 324 
    -- successors 326 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__condition_check__/$exit
      -- 
    cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(318) & cp_elements(324);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(325), clk => clk, reset => reset); --
    end block;
    Xexit_9722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => switch_stmt_2045_branch_default_req_0); -- 
    -- CP-element group 326 branch  place  bypass 
    -- predecessors 325 
    -- successors 327 329 331 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045__select__
      -- 
    cp_elements(326) <= cp_elements(325);
    -- CP-element group 327 transition  bypass 
    -- predecessors 326 
    -- successors 328 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_0/$entry
      -- 
    cp_elements(327) <= cp_elements(326);
    -- CP-element group 328 fork  transition  place  input  bypass 
    -- predecessors 327 
    -- successors 1400 1401 
    -- members (8) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_0/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_0/ack1
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/$entry
      -- 
    ack1_9761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_branch_0_ack_1, ack => cp_elements(328)); -- 
    -- CP-element group 329 transition  bypass 
    -- predecessors 326 
    -- successors 330 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_1/$entry
      -- 
    cp_elements(329) <= cp_elements(326);
    -- CP-element group 330 fork  transition  place  input  bypass 
    -- predecessors 329 
    -- successors 1411 1415 
    -- members (6) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_1/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_1/ack1
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- 
    ack1_9766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_branch_1_ack_1, ack => cp_elements(330)); -- 
    -- CP-element group 331 transition  bypass 
    -- predecessors 326 
    -- successors 332 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_default/$entry
      -- 
    cp_elements(331) <= cp_elements(326);
    -- CP-element group 332 transition  place  input  bypass 
    -- predecessors 331 
    -- successors 12 
    -- members (9) 
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_default/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2045_choice_default/ack0
      -- 	branch_block_stmt_1659/bb_12_bbx_xnph7x_xix_xix_xi5x_xpreheader
      -- 	branch_block_stmt_1659/bb_12_bbx_xnph7x_xix_xix_xi5x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_12_bbx_xnph7x_xix_xix_xi5x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2055_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_2055_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2055_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2055_PhiAck/dummy
      -- 
    ack0_9771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2045_branch_default_ack_0, ack => cp_elements(332)); -- 
    -- CP-element group 333 fork  transition  bypass 
    -- predecessors 13 
    -- successors 334 335 339 340 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/$entry
      -- 
    cp_elements(333) <= cp_elements(13);
    -- CP-element group 334 transition  output  bypass 
    -- predecessors 333 
    -- successors 337 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Update/cr
      -- 
    cp_elements(334) <= cp_elements(333);
    cr_9792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(334), ack => LSHR_u32_u32_2076_inst_req_1); -- 
    -- CP-element group 335 transition  output  bypass 
    -- predecessors 333 
    -- successors 336 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_xx_x016x_xix_xix_xi3_2073_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_xx_x016x_xix_xix_xi3_2073_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_xx_x016x_xix_xix_xi3_2073_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_xx_x016x_xix_xix_xi3_2073_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Sample/rr
      -- 
    cp_elements(335) <= cp_elements(333);
    rr_9787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => LSHR_u32_u32_2076_inst_req_0); -- 
    -- CP-element group 336 transition  input  bypass 
    -- predecessors 335 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Sample/ra
      -- 
    ra_9788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2076_inst_ack_0, ack => cp_elements(336)); -- 
    -- CP-element group 337 transition  input  bypass 
    -- predecessors 334 
    -- successors 338 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/LSHR_u32_u32_2076_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_108_2079_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_108_2079_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_108_2079_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_108_2079_update_completed_
      -- 
    ca_9793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2076_inst_ack_1, ack => cp_elements(337)); -- 
    -- CP-element group 338 join  transition  output  bypass 
    -- predecessors 337 340 
    -- successors 341 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Sample/rr
      -- 
    cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(337) & cp_elements(340);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(338), clk => clk, reset => reset); --
    end block;
    rr_9809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => UGT_u32_u1_2081_inst_req_0); -- 
    -- CP-element group 339 transition  output  bypass 
    -- predecessors 333 
    -- successors 342 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Update/cr
      -- 
    cp_elements(339) <= cp_elements(333);
    cr_9814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => UGT_u32_u1_2081_inst_req_1); -- 
    -- CP-element group 340 transition  bypass 
    -- predecessors 333 
    -- successors 338 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_61_2080_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_61_2080_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_61_2080_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/R_iNsTr_61_2080_update_completed_
      -- 
    cp_elements(340) <= cp_elements(333);
    -- CP-element group 341 transition  input  bypass 
    -- predecessors 338 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Sample/ra
      -- 
    ra_9810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2081_inst_ack_0, ack => cp_elements(341)); -- 
    -- CP-element group 342 branch  transition  place  input  bypass 
    -- predecessors 339 
    -- successors 343 344 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2083__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2077_to_assign_stmt_2082/UGT_u32_u1_2081_Update/ca
      -- 
    ca_9815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2081_inst_ack_1, ack => cp_elements(342)); -- 
    -- CP-element group 343 transition  place  dead  bypass 
    -- predecessors 342 
    -- successors 14 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2083__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2089__entry__
      -- 	branch_block_stmt_1659/if_stmt_2083_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2083_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2083_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2089_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2089_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2089_dead_link/dead_transition
      -- 
    cp_elements(343) <= false;
    -- CP-element group 344 transition  output  bypass 
    -- predecessors 342 
    -- successors 345 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2083_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2083_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2083_eval_test/branch_req
      -- 
    cp_elements(344) <= cp_elements(342);
    branch_req_9823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(344), ack => if_stmt_2083_branch_req_0); -- 
    -- CP-element group 345 branch  place  bypass 
    -- predecessors 344 
    -- successors 346 348 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_109_2084_place
      -- 
    cp_elements(345) <= cp_elements(344);
    -- CP-element group 346 transition  bypass 
    -- predecessors 345 
    -- successors 347 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2083_if_link/$entry
      -- 
    cp_elements(346) <= cp_elements(345);
    -- CP-element group 347 transition  place  input  bypass 
    -- predecessors 346 
    -- successors 14 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2083_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2083_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_bbx_xnphx_xix_xix_xi8x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2089_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_2089_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2089_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2089_PhiAck/dummy
      -- 
    if_choice_transition_9828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2083_branch_ack_1, ack => cp_elements(347)); -- 
    -- CP-element group 348 transition  bypass 
    -- predecessors 345 
    -- successors 349 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2083_else_link/$entry
      -- 
    cp_elements(348) <= cp_elements(345);
    -- CP-element group 349 transition  place  input  bypass 
    -- predecessors 348 
    -- successors 1351 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2083_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2083_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11
      -- 
    else_choice_transition_9832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2083_branch_ack_0, ack => cp_elements(349)); -- 
    -- CP-element group 350 fork  transition  bypass 
    -- predecessors 15 
    -- successors 351 352 355 356 360 361 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/$entry
      -- 
    cp_elements(350) <= cp_elements(15);
    -- CP-element group 351 transition  output  bypass 
    -- predecessors 350 
    -- successors 354 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Update/cr
      -- 
    cp_elements(351) <= cp_elements(350);
    cr_9854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => SHL_u32_u32_2110_inst_req_1); -- 
    -- CP-element group 352 transition  output  bypass 
    -- predecessors 350 
    -- successors 353 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_shifted_divisorx_x03x_xix_xix_xi6_2107_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_shifted_divisorx_x03x_xix_xix_xi6_2107_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_shifted_divisorx_x03x_xix_xix_xi6_2107_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_shifted_divisorx_x03x_xix_xix_xi6_2107_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Sample/rr
      -- 
    cp_elements(352) <= cp_elements(350);
    rr_9849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(352), ack => SHL_u32_u32_2110_inst_req_0); -- 
    -- CP-element group 353 transition  input  bypass 
    -- predecessors 352 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Sample/ra
      -- 
    ra_9850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2110_inst_ack_0, ack => cp_elements(353)); -- 
    -- CP-element group 354 transition  input  bypass 
    -- predecessors 351 
    -- successors 359 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2110_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_162_2119_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_162_2119_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_162_2119_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_162_2119_update_completed_
      -- 
    ca_9855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2110_inst_ack_1, ack => cp_elements(354)); -- 
    -- CP-element group 355 transition  output  bypass 
    -- predecessors 350 
    -- successors 358 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Update/cr
      -- 
    cp_elements(355) <= cp_elements(350);
    cr_9872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(355), ack => SHL_u32_u32_2116_inst_req_1); -- 
    -- CP-element group 356 transition  output  bypass 
    -- predecessors 350 
    -- successors 357 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_curr_quotientx_x02x_xix_xix_xi7_2113_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_curr_quotientx_x02x_xix_xix_xi7_2113_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_curr_quotientx_x02x_xix_xix_xi7_2113_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_curr_quotientx_x02x_xix_xix_xi7_2113_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Sample/rr
      -- 
    cp_elements(356) <= cp_elements(350);
    rr_9867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => SHL_u32_u32_2116_inst_req_0); -- 
    -- CP-element group 357 transition  input  bypass 
    -- predecessors 356 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Sample/ra
      -- 
    ra_9868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2116_inst_ack_0, ack => cp_elements(357)); -- 
    -- CP-element group 358 transition  input  bypass 
    -- predecessors 355 
    -- successors 364 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/SHL_u32_u32_2116_Update/ca
      -- 
    ca_9873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2116_inst_ack_1, ack => cp_elements(358)); -- 
    -- CP-element group 359 join  transition  output  bypass 
    -- predecessors 354 361 
    -- successors 362 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Sample/rr
      -- 
    cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(354) & cp_elements(361);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(359), clk => clk, reset => reset); --
    end block;
    rr_9889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(359), ack => ULT_u32_u1_2121_inst_req_0); -- 
    -- CP-element group 360 transition  output  bypass 
    -- predecessors 350 
    -- successors 363 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Update/cr
      -- 
    cp_elements(360) <= cp_elements(350);
    cr_9894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => ULT_u32_u1_2121_inst_req_1); -- 
    -- CP-element group 361 transition  bypass 
    -- predecessors 350 
    -- successors 359 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_108_2120_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_108_2120_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_108_2120_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/R_iNsTr_108_2120_update_completed_
      -- 
    cp_elements(361) <= cp_elements(350);
    -- CP-element group 362 transition  input  bypass 
    -- predecessors 359 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Sample/ra
      -- 
    ra_9890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2121_inst_ack_0, ack => cp_elements(362)); -- 
    -- CP-element group 363 transition  input  bypass 
    -- predecessors 360 
    -- successors 364 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/ULT_u32_u1_2121_Update/ca
      -- 
    ca_9895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2121_inst_ack_1, ack => cp_elements(363)); -- 
    -- CP-element group 364 join  transition  bypass 
    -- predecessors 358 363 
    -- successors 16 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2111_to_assign_stmt_2122/$exit
      -- 
    cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(358) & cp_elements(363);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365 transition  place  dead  bypass 
    -- predecessors 16 
    -- successors 17 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2129__entry__
      -- 	branch_block_stmt_1659/if_stmt_2123__exit__
      -- 	branch_block_stmt_1659/if_stmt_2123_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2123_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2123_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2129_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2129_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2129_dead_link/dead_transition
      -- 
    cp_elements(365) <= false;
    -- CP-element group 366 transition  output  bypass 
    -- predecessors 16 
    -- successors 367 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2123_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2123_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2123_eval_test/branch_req
      -- 
    cp_elements(366) <= cp_elements(16);
    branch_req_9903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(366), ack => if_stmt_2123_branch_req_0); -- 
    -- CP-element group 367 branch  place  bypass 
    -- predecessors 366 
    -- successors 368 370 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_164_2124_place
      -- 
    cp_elements(367) <= cp_elements(366);
    -- CP-element group 368 transition  bypass 
    -- predecessors 367 
    -- successors 369 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2123_if_link/$entry
      -- 
    cp_elements(368) <= cp_elements(367);
    -- CP-element group 369 transition  place  input  bypass 
    -- predecessors 368 
    -- successors 1289 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2123_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2123_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8
      -- 
    if_choice_transition_9908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2123_branch_ack_1, ack => cp_elements(369)); -- 
    -- CP-element group 370 transition  bypass 
    -- predecessors 367 
    -- successors 371 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2123_else_link/$entry
      -- 
    cp_elements(370) <= cp_elements(367);
    -- CP-element group 371 transition  place  input  bypass 
    -- predecessors 370 
    -- successors 1332 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2123_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2123_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit
      -- 
    else_choice_transition_9912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2123_branch_ack_0, ack => cp_elements(371)); -- 
    -- CP-element group 372 fork  transition  bypass 
    -- predecessors 18 
    -- successors 374 375 376 380 381 382 386 387 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/$entry
      -- 
    cp_elements(372) <= cp_elements(18);
    -- CP-element group 373 join  transition  output  bypass 
    -- predecessors 375 376 
    -- successors 377 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Sample/rr
      -- 
    cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(375) & cp_elements(376);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(373), clk => clk, reset => reset); --
    end block;
    rr_9933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(373), ack => ADD_u32_u32_2158_inst_req_0); -- 
    -- CP-element group 374 transition  output  bypass 
    -- predecessors 372 
    -- successors 378 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Update/cr
      -- 
    cp_elements(374) <= cp_elements(372);
    cr_9938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(374), ack => ADD_u32_u32_2158_inst_req_1); -- 
    -- CP-element group 375 transition  bypass 
    -- predecessors 372 
    -- successors 373 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2156_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2156_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2156_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_curr_quotientx_x0x_xlcssax_xix_xix_xi10_2156_update_completed_
      -- 
    cp_elements(375) <= cp_elements(372);
    -- CP-element group 376 transition  bypass 
    -- predecessors 372 
    -- successors 373 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_quotientx_x05x_xix_xix_xi4_2157_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_quotientx_x05x_xix_xix_xi4_2157_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_quotientx_x05x_xix_xix_xi4_2157_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_quotientx_x05x_xix_xix_xi4_2157_update_completed_
      -- 
    cp_elements(376) <= cp_elements(372);
    -- CP-element group 377 transition  input  bypass 
    -- predecessors 373 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Sample/ra
      -- 
    ra_9934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2158_inst_ack_0, ack => cp_elements(377)); -- 
    -- CP-element group 378 transition  input  bypass 
    -- predecessors 374 
    -- successors 390 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ADD_u32_u32_2158_Update/ca
      -- 
    ca_9939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2158_inst_ack_1, ack => cp_elements(378)); -- 
    -- CP-element group 379 join  transition  output  bypass 
    -- predecessors 381 382 
    -- successors 383 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Sample/rr
      -- 
    cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(381) & cp_elements(382);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(379), clk => clk, reset => reset); --
    end block;
    rr_9955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => SUB_u32_u32_2163_inst_req_0); -- 
    -- CP-element group 380 transition  output  bypass 
    -- predecessors 372 
    -- successors 384 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Update/cr
      -- 
    cp_elements(380) <= cp_elements(372);
    cr_9960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => SUB_u32_u32_2163_inst_req_1); -- 
    -- CP-element group 381 transition  bypass 
    -- predecessors 372 
    -- successors 379 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_xx_x016x_xix_xix_xi3_2161_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_xx_x016x_xix_xix_xi3_2161_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_xx_x016x_xix_xix_xi3_2161_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_xx_x016x_xix_xix_xi3_2161_update_completed_
      -- 
    cp_elements(381) <= cp_elements(372);
    -- CP-element group 382 transition  bypass 
    -- predecessors 372 
    -- successors 379 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2162_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2162_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2162_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2162_update_completed_
      -- 
    cp_elements(382) <= cp_elements(372);
    -- CP-element group 383 transition  input  bypass 
    -- predecessors 379 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Sample/ra
      -- 
    ra_9956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2163_inst_ack_0, ack => cp_elements(383)); -- 
    -- CP-element group 384 transition  input  bypass 
    -- predecessors 380 
    -- successors 385 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/SUB_u32_u32_2163_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_137_2166_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_137_2166_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_137_2166_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_137_2166_update_completed_
      -- 
    ca_9961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2163_inst_ack_1, ack => cp_elements(384)); -- 
    -- CP-element group 385 join  transition  output  bypass 
    -- predecessors 384 387 
    -- successors 388 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Sample/rr
      -- 
    cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(384) & cp_elements(387);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(385), clk => clk, reset => reset); --
    end block;
    rr_9977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(385), ack => ULT_u32_u1_2168_inst_req_0); -- 
    -- CP-element group 386 transition  output  bypass 
    -- predecessors 372 
    -- successors 389 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Update/cr
      -- 
    cp_elements(386) <= cp_elements(372);
    cr_9982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => ULT_u32_u1_2168_inst_req_1); -- 
    -- CP-element group 387 transition  bypass 
    -- predecessors 372 
    -- successors 385 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_61_2167_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_61_2167_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_61_2167_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/R_iNsTr_61_2167_update_completed_
      -- 
    cp_elements(387) <= cp_elements(372);
    -- CP-element group 388 transition  input  bypass 
    -- predecessors 385 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Sample/ra
      -- 
    ra_9978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2168_inst_ack_0, ack => cp_elements(388)); -- 
    -- CP-element group 389 transition  input  bypass 
    -- predecessors 386 
    -- successors 390 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/ULT_u32_u1_2168_Update/ca
      -- 
    ca_9983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2168_inst_ack_1, ack => cp_elements(389)); -- 
    -- CP-element group 390 join  transition  bypass 
    -- predecessors 378 389 
    -- successors 19 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2159_to_assign_stmt_2169/$exit
      -- 
    cp_element_group_390: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_390"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(378) & cp_elements(389);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(390), clk => clk, reset => reset); --
    end block;
    -- CP-element group 391 transition  place  dead  bypass 
    -- predecessors 19 
    -- successors 20 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2170__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2176__entry__
      -- 	branch_block_stmt_1659/if_stmt_2170_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2170_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2170_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2176_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2176_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2176_dead_link/$entry
      -- 
    cp_elements(391) <= false;
    -- CP-element group 392 transition  output  bypass 
    -- predecessors 19 
    -- successors 393 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2170_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2170_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2170_eval_test/branch_req
      -- 
    cp_elements(392) <= cp_elements(19);
    branch_req_9991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(392), ack => if_stmt_2170_branch_req_0); -- 
    -- CP-element group 393 branch  place  bypass 
    -- predecessors 392 
    -- successors 394 396 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_138_2171_place
      -- 
    cp_elements(393) <= cp_elements(392);
    -- CP-element group 394 transition  bypass 
    -- predecessors 393 
    -- successors 395 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2170_if_link/$entry
      -- 
    cp_elements(394) <= cp_elements(393);
    -- CP-element group 395 fork  transition  place  input  bypass 
    -- predecessors 394 
    -- successors 1394 1396 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2170_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2170_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_9996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2170_branch_ack_1, ack => cp_elements(395)); -- 
    -- CP-element group 396 transition  bypass 
    -- predecessors 393 
    -- successors 397 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2170_else_link/$entry
      -- 
    cp_elements(396) <= cp_elements(393);
    -- CP-element group 397 transition  place  input  bypass 
    -- predecessors 396 
    -- successors 1264 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2170_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2170_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5
      -- 
    else_choice_transition_10000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2170_branch_ack_0, ack => cp_elements(397)); -- 
    -- CP-element group 398 fork  transition  bypass 
    -- predecessors 1435 
    -- successors 399 400 403 406 407 413 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/$entry
      -- 
    cp_elements(398) <= cp_elements(1435);
    -- CP-element group 399 transition  output  bypass 
    -- predecessors 398 
    -- successors 402 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Update/cr
      -- 
    cp_elements(399) <= cp_elements(398);
    cr_10022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(399), ack => AND_u32_u32_2205_inst_req_1); -- 
    -- CP-element group 400 transition  output  bypass 
    -- predecessors 398 
    -- successors 401 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2202_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2202_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2202_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2202_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Sample/rr
      -- 
    cp_elements(400) <= cp_elements(398);
    rr_10017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => AND_u32_u32_2205_inst_req_0); -- 
    -- CP-element group 401 transition  input  bypass 
    -- predecessors 400 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Sample/ra
      -- 
    ra_10018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2205_inst_ack_0, ack => cp_elements(401)); -- 
    -- CP-element group 402 transition  input  output  bypass 
    -- predecessors 399 
    -- successors 404 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u32_u32_2205_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_92_2208_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_92_2208_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_92_2208_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_92_2208_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Sample/rr
      -- 
    ca_10023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2205_inst_ack_1, ack => cp_elements(402)); -- 
    rr_10035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => EQ_u32_u1_2211_inst_req_0); -- 
    -- CP-element group 403 transition  output  bypass 
    -- predecessors 398 
    -- successors 405 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Update/cr
      -- 
    cp_elements(403) <= cp_elements(398);
    cr_10040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(403), ack => EQ_u32_u1_2211_inst_req_1); -- 
    -- CP-element group 404 transition  input  bypass 
    -- predecessors 402 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Sample/ra
      -- 
    ra_10036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2211_inst_ack_0, ack => cp_elements(404)); -- 
    -- CP-element group 405 transition  input  bypass 
    -- predecessors 403 
    -- successors 412 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/EQ_u32_u1_2211_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_93_2222_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_93_2222_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_93_2222_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_93_2222_update_completed_
      -- 
    ca_10041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2211_inst_ack_1, ack => cp_elements(405)); -- 
    -- CP-element group 406 transition  output  bypass 
    -- predecessors 398 
    -- successors 411 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Update/cr
      -- 
    cp_elements(406) <= cp_elements(398);
    cr_10072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => NEQ_i32_u1_2219_inst_req_1); -- 
    -- CP-element group 407 transition  output  bypass 
    -- predecessors 398 
    -- successors 408 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2214_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2214_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2214_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_tempx_x0x_xphx_xix_xi14_2214_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Sample/rr
      -- 
    cp_elements(407) <= cp_elements(398);
    rr_10057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => type_cast_2215_inst_req_0); -- 
    -- CP-element group 408 transition  input  output  bypass 
    -- predecessors 407 
    -- successors 409 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Update/cr
      -- 
    ra_10058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_0, ack => cp_elements(408)); -- 
    cr_10062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(408), ack => type_cast_2215_inst_req_1); -- 
    -- CP-element group 409 transition  input  output  bypass 
    -- predecessors 408 
    -- successors 410 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/type_cast_2215_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Sample/rr
      -- 
    ca_10063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_1, ack => cp_elements(409)); -- 
    rr_10067_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(409), ack => NEQ_i32_u1_2219_inst_req_0); -- 
    -- CP-element group 410 transition  input  bypass 
    -- predecessors 409 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Sample/ra
      -- 
    ra_10068_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2219_inst_ack_0, ack => cp_elements(410)); -- 
    -- CP-element group 411 transition  input  bypass 
    -- predecessors 406 
    -- successors 412 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/NEQ_i32_u1_2219_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_94_2223_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_94_2223_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_94_2223_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/R_iNsTr_94_2223_update_completed_
      -- 
    ca_10073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2219_inst_ack_1, ack => cp_elements(411)); -- 
    -- CP-element group 412 join  transition  output  bypass 
    -- predecessors 405 411 
    -- successors 414 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Sample/rr
      -- 
    cp_element_group_412: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_412"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(405) & cp_elements(411);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(412), clk => clk, reset => reset); --
    end block;
    rr_10089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(412), ack => AND_u1_u1_2224_inst_req_0); -- 
    -- CP-element group 413 transition  output  bypass 
    -- predecessors 398 
    -- successors 415 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Update/cr
      -- 
    cp_elements(413) <= cp_elements(398);
    cr_10094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(413), ack => AND_u1_u1_2224_inst_req_1); -- 
    -- CP-element group 414 transition  input  bypass 
    -- predecessors 412 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Sample/ra
      -- 
    ra_10090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2224_inst_ack_0, ack => cp_elements(414)); -- 
    -- CP-element group 415 branch  transition  place  input  bypass 
    -- predecessors 413 
    -- successors 416 417 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2226__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225/AND_u1_u1_2224_Update/ca
      -- 
    ca_10095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2224_inst_ack_1, ack => cp_elements(415)); -- 
    -- CP-element group 416 transition  place  dead  bypass 
    -- predecessors 415 
    -- successors 21 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2232__entry__
      -- 	branch_block_stmt_1659/if_stmt_2226__exit__
      -- 	branch_block_stmt_1659/if_stmt_2226_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2226_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2226_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2232_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2232_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2232_dead_link/dead_transition
      -- 
    cp_elements(416) <= false;
    -- CP-element group 417 transition  output  bypass 
    -- predecessors 415 
    -- successors 418 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2226_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2226_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2226_eval_test/branch_req
      -- 
    cp_elements(417) <= cp_elements(415);
    branch_req_10103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(417), ack => if_stmt_2226_branch_req_0); -- 
    -- CP-element group 418 branch  place  bypass 
    -- predecessors 417 
    -- successors 419 421 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcond11x_xix_xi15_2227_place
      -- 
    cp_elements(418) <= cp_elements(417);
    -- CP-element group 419 transition  bypass 
    -- predecessors 418 
    -- successors 420 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2226_if_link/$entry
      -- 
    cp_elements(419) <= cp_elements(418);
    -- CP-element group 420 transition  place  input  bypass 
    -- predecessors 419 
    -- successors 21 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2226_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2226_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader
      -- 	branch_block_stmt_1659/merge_stmt_2232_PhiReqMerge
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_udiv32x_xexitx_xix_xi20x_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2232_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2232_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2232_PhiAck/dummy
      -- 
    if_choice_transition_10108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2226_branch_ack_1, ack => cp_elements(420)); -- 
    -- CP-element group 421 transition  bypass 
    -- predecessors 418 
    -- successors 422 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2226_else_link/$entry
      -- 
    cp_elements(421) <= cp_elements(418);
    -- CP-element group 422 transition  place  input  bypass 
    -- predecessors 421 
    -- successors 1498 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2226_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2226_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29
      -- 
    else_choice_transition_10112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2226_branch_ack_0, ack => cp_elements(422)); -- 
    -- CP-element group 423 fork  transition  bypass 
    -- predecessors 22 
    -- successors 424 425 428 432 435 442 445 446 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/$entry
      -- 
    cp_elements(423) <= cp_elements(22);
    -- CP-element group 424 transition  output  bypass 
    -- predecessors 423 
    -- successors 427 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Update/cr
      -- 
    cp_elements(424) <= cp_elements(423);
    cr_10134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(424), ack => SHL_u32_u32_2253_inst_req_1); -- 
    -- CP-element group 425 transition  output  bypass 
    -- predecessors 423 
    -- successors 426 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_tempx_x012x_xix_xi17_2250_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_tempx_x012x_xix_xi17_2250_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_tempx_x012x_xix_xi17_2250_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_tempx_x012x_xix_xi17_2250_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Sample/rr
      -- 
    cp_elements(425) <= cp_elements(423);
    rr_10129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(425), ack => SHL_u32_u32_2253_inst_req_0); -- 
    -- CP-element group 426 transition  input  bypass 
    -- predecessors 425 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Sample/ra
      -- 
    ra_10130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2253_inst_ack_0, ack => cp_elements(426)); -- 
    -- CP-element group 427 fork  transition  input  bypass 
    -- predecessors 424 
    -- successors 429 436 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/SHL_u32_u32_2253_Update/ca
      -- 
    ca_10135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2253_inst_ack_1, ack => cp_elements(427)); -- 
    -- CP-element group 428 transition  output  bypass 
    -- predecessors 423 
    -- successors 431 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Update/cr
      -- 
    cp_elements(428) <= cp_elements(423);
    cr_10152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => AND_u32_u32_2259_inst_req_1); -- 
    -- CP-element group 429 transition  output  bypass 
    -- predecessors 427 
    -- successors 430 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2256_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2256_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2256_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2256_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Sample/rr
      -- 
    cp_elements(429) <= cp_elements(427);
    rr_10147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(429), ack => AND_u32_u32_2259_inst_req_0); -- 
    -- CP-element group 430 transition  input  bypass 
    -- predecessors 429 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Sample/ra
      -- 
    ra_10148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2259_inst_ack_0, ack => cp_elements(430)); -- 
    -- CP-element group 431 transition  input  output  bypass 
    -- predecessors 428 
    -- successors 433 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u32_u32_2259_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_142_2262_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_142_2262_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_142_2262_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_142_2262_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Sample/rr
      -- 
    ca_10153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2259_inst_ack_1, ack => cp_elements(431)); -- 
    rr_10165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(431), ack => EQ_u32_u1_2265_inst_req_0); -- 
    -- CP-element group 432 transition  output  bypass 
    -- predecessors 423 
    -- successors 434 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Update/cr
      -- 
    cp_elements(432) <= cp_elements(423);
    cr_10170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(432), ack => EQ_u32_u1_2265_inst_req_1); -- 
    -- CP-element group 433 transition  input  bypass 
    -- predecessors 431 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Sample/ra
      -- 
    ra_10166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2265_inst_ack_0, ack => cp_elements(433)); -- 
    -- CP-element group 434 transition  input  bypass 
    -- predecessors 432 
    -- successors 441 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/EQ_u32_u1_2265_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_143_2276_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_143_2276_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_143_2276_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_143_2276_update_completed_
      -- 
    ca_10171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2265_inst_ack_1, ack => cp_elements(434)); -- 
    -- CP-element group 435 transition  output  bypass 
    -- predecessors 423 
    -- successors 440 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Update/cr
      -- 
    cp_elements(435) <= cp_elements(423);
    cr_10202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => NEQ_i32_u1_2273_inst_req_1); -- 
    -- CP-element group 436 transition  output  bypass 
    -- predecessors 427 
    -- successors 437 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2268_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2268_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2268_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_141_2268_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Sample/rr
      -- 
    cp_elements(436) <= cp_elements(427);
    rr_10187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => type_cast_2269_inst_req_0); -- 
    -- CP-element group 437 transition  input  output  bypass 
    -- predecessors 436 
    -- successors 438 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Update/cr
      -- 
    ra_10188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_0, ack => cp_elements(437)); -- 
    cr_10192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(437), ack => type_cast_2269_inst_req_1); -- 
    -- CP-element group 438 transition  input  output  bypass 
    -- predecessors 437 
    -- successors 439 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/type_cast_2269_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Sample/rr
      -- 
    ca_10193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_1, ack => cp_elements(438)); -- 
    rr_10197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => NEQ_i32_u1_2273_inst_req_0); -- 
    -- CP-element group 439 transition  input  bypass 
    -- predecessors 438 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Sample/ra
      -- 
    ra_10198_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2273_inst_ack_0, ack => cp_elements(439)); -- 
    -- CP-element group 440 transition  input  bypass 
    -- predecessors 435 
    -- successors 441 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/NEQ_i32_u1_2273_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_144_2277_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_144_2277_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_144_2277_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_144_2277_update_completed_
      -- 
    ca_10203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2273_inst_ack_1, ack => cp_elements(440)); -- 
    -- CP-element group 441 join  transition  output  bypass 
    -- predecessors 434 440 
    -- successors 443 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Sample/rr
      -- 
    cp_element_group_441: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_441"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(434) & cp_elements(440);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(441), clk => clk, reset => reset); --
    end block;
    rr_10219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => AND_u1_u1_2278_inst_req_0); -- 
    -- CP-element group 442 transition  output  bypass 
    -- predecessors 423 
    -- successors 444 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Update/cr
      -- 
    cp_elements(442) <= cp_elements(423);
    cr_10224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => AND_u1_u1_2278_inst_req_1); -- 
    -- CP-element group 443 transition  input  bypass 
    -- predecessors 441 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Sample/ra
      -- 
    ra_10220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2278_inst_ack_0, ack => cp_elements(443)); -- 
    -- CP-element group 444 transition  input  bypass 
    -- predecessors 442 
    -- successors 449 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/AND_u1_u1_2278_Update/ca
      -- 
    ca_10225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2278_inst_ack_1, ack => cp_elements(444)); -- 
    -- CP-element group 445 transition  output  bypass 
    -- predecessors 423 
    -- successors 448 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_update_start_
      -- 
    cp_elements(445) <= cp_elements(423);
    cr_10242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => ADD_u32_u32_2284_inst_req_1); -- 
    -- CP-element group 446 transition  output  bypass 
    -- predecessors 423 
    -- successors 447 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_140_2281_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_140_2281_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_140_2281_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/R_iNsTr_140_2281_sample_start_
      -- 
    cp_elements(446) <= cp_elements(423);
    rr_10237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(446), ack => ADD_u32_u32_2284_inst_req_0); -- 
    -- CP-element group 447 transition  input  bypass 
    -- predecessors 446 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_sample_completed_
      -- 
    ra_10238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2284_inst_ack_0, ack => cp_elements(447)); -- 
    -- CP-element group 448 transition  input  bypass 
    -- predecessors 445 
    -- successors 449 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/ADD_u32_u32_2284_update_completed_
      -- 
    ca_10243_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2284_inst_ack_1, ack => cp_elements(448)); -- 
    -- CP-element group 449 join  transition  bypass 
    -- predecessors 444 448 
    -- successors 23 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2254_to_assign_stmt_2285/$exit
      -- 
    cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(444) & cp_elements(448);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450 transition  place  dead  bypass 
    -- predecessors 23 
    -- successors 24 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2286__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2292__entry__
      -- 	branch_block_stmt_1659/if_stmt_2286_dead_link/dead_transition
      -- 	branch_block_stmt_1659/if_stmt_2286_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2286_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2292_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2292_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2292_dead_link/dead_transition
      -- 
    cp_elements(450) <= false;
    -- CP-element group 451 transition  output  bypass 
    -- predecessors 23 
    -- successors 452 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2286_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2286_eval_test/branch_req
      -- 	branch_block_stmt_1659/if_stmt_2286_eval_test/$exit
      -- 
    cp_elements(451) <= cp_elements(23);
    branch_req_10251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(451), ack => if_stmt_2286_branch_req_0); -- 
    -- CP-element group 452 branch  place  bypass 
    -- predecessors 451 
    -- successors 453 455 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcondx_xix_xi18_2287_place
      -- 
    cp_elements(452) <= cp_elements(451);
    -- CP-element group 453 transition  bypass 
    -- predecessors 452 
    -- successors 454 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2286_if_link/$entry
      -- 
    cp_elements(453) <= cp_elements(452);
    -- CP-element group 454 transition  place  input  bypass 
    -- predecessors 453 
    -- successors 1436 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2286_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/if_stmt_2286_if_link/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20
      -- 
    if_choice_transition_10256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2286_branch_ack_1, ack => cp_elements(454)); -- 
    -- CP-element group 455 transition  bypass 
    -- predecessors 452 
    -- successors 456 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2286_else_link/$entry
      -- 
    cp_elements(455) <= cp_elements(452);
    -- CP-element group 456 transition  place  input  bypass 
    -- predecessors 455 
    -- successors 1479 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25
      -- 	branch_block_stmt_1659/if_stmt_2286_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/if_stmt_2286_else_link/$exit
      -- 
    else_choice_transition_10260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2286_branch_ack_0, ack => cp_elements(456)); -- 
    -- CP-element group 457 fork  transition  bypass 
    -- predecessors 24 
    -- successors 458 459 462 466 467 471 472 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/$entry
      -- 
    cp_elements(457) <= cp_elements(24);
    -- CP-element group 458 transition  output  bypass 
    -- predecessors 457 
    -- successors 461 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_update_start_
      -- 
    cp_elements(458) <= cp_elements(457);
    cr_10282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => OR_u32_u32_2306_inst_req_1); -- 
    -- CP-element group 459 transition  output  bypass 
    -- predecessors 457 
    -- successors 460 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_54_2303_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_54_2303_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_54_2303_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_54_2303_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_sample_start_
      -- 
    cp_elements(459) <= cp_elements(457);
    rr_10277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(459), ack => OR_u32_u32_2306_inst_req_0); -- 
    -- CP-element group 460 transition  input  bypass 
    -- predecessors 459 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_sample_completed_
      -- 
    ra_10278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2306_inst_ack_0, ack => cp_elements(460)); -- 
    -- CP-element group 461 transition  input  output  bypass 
    -- predecessors 458 
    -- successors 463 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xnotx_xi21_2309_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xnotx_xi21_2309_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xnotx_xi21_2309_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xnotx_xi21_2309_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/OR_u32_u32_2306_update_completed_
      -- 
    ca_10283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2306_inst_ack_1, ack => cp_elements(461)); -- 
    rr_10295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => XOR_u32_u32_2312_inst_req_0); -- 
    -- CP-element group 462 transition  output  bypass 
    -- predecessors 457 
    -- successors 464 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_update_start_
      -- 
    cp_elements(462) <= cp_elements(457);
    cr_10300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => XOR_u32_u32_2312_inst_req_1); -- 
    -- CP-element group 463 transition  input  bypass 
    -- predecessors 461 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_sample_completed_
      -- 
    ra_10296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2312_inst_ack_0, ack => cp_elements(463)); -- 
    -- CP-element group 464 transition  input  bypass 
    -- predecessors 462 
    -- successors 465 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp21x_xix_xi22_2315_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp21x_xix_xi22_2315_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp21x_xix_xi22_2315_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp21x_xix_xi22_2315_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/XOR_u32_u32_2312_update_completed_
      -- 
    ca_10301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2312_inst_ack_1, ack => cp_elements(464)); -- 
    -- CP-element group 465 join  transition  output  bypass 
    -- predecessors 464 467 
    -- successors 468 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Sample/rr
      -- 
    cp_element_group_465: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_465"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(464) & cp_elements(467);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(465), clk => clk, reset => reset); --
    end block;
    rr_10317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(465), ack => ADD_u32_u32_2317_inst_req_0); -- 
    -- CP-element group 466 transition  output  bypass 
    -- predecessors 457 
    -- successors 469 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Update/$entry
      -- 
    cp_elements(466) <= cp_elements(457);
    cr_10322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => ADD_u32_u32_2317_inst_req_1); -- 
    -- CP-element group 467 transition  bypass 
    -- predecessors 457 
    -- successors 465 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_53_2316_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_53_2316_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_53_2316_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_iNsTr_53_2316_update_start_
      -- 
    cp_elements(467) <= cp_elements(457);
    -- CP-element group 468 transition  input  bypass 
    -- predecessors 465 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Sample/$exit
      -- 
    ra_10318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2317_inst_ack_0, ack => cp_elements(468)); -- 
    -- CP-element group 469 transition  input  bypass 
    -- predecessors 466 
    -- successors 470 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp25x_xix_xi23_2320_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp25x_xix_xi23_2320_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp25x_xix_xi23_2320_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/ADD_u32_u32_2317_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_tmp25x_xix_xi23_2320_sample_completed_
      -- 
    ca_10323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2317_inst_ack_1, ack => cp_elements(469)); -- 
    -- CP-element group 470 join  transition  output  bypass 
    -- predecessors 469 472 
    -- successors 473 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Sample/$entry
      -- 
    cp_element_group_470: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_470"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(469) & cp_elements(472);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(470), clk => clk, reset => reset); --
    end block;
    rr_10339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(470), ack => SUB_u32_u32_2322_inst_req_0); -- 
    -- CP-element group 471 transition  output  bypass 
    -- predecessors 457 
    -- successors 474 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Update/cr
      -- 
    cp_elements(471) <= cp_elements(457);
    cr_10344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(471), ack => SUB_u32_u32_2322_inst_req_1); -- 
    -- CP-element group 472 transition  bypass 
    -- predecessors 457 
    -- successors 470 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xlcssa10_2321_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xlcssa10_2321_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xlcssa10_2321_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/R_xx_xlcssa10_2321_update_completed_
      -- 
    cp_elements(472) <= cp_elements(457);
    -- CP-element group 473 transition  input  bypass 
    -- predecessors 470 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Sample/$exit
      -- 
    ra_10340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2322_inst_ack_0, ack => cp_elements(473)); -- 
    -- CP-element group 474 transition  place  input  bypass 
    -- predecessors 471 
    -- successors 1524 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323__exit__
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2307_to_assign_stmt_2323/SUB_u32_u32_2322_Update/ca
      -- 
    ca_10345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2322_inst_ack_1, ack => cp_elements(474)); -- 
    -- CP-element group 475 fork  transition  bypass 
    -- predecessors 25 
    -- successors 476 477 480 481 484 488 489 493 496 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/$entry
      -- 
    cp_elements(475) <= cp_elements(25);
    -- CP-element group 476 transition  output  bypass 
    -- predecessors 475 
    -- successors 479 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Update/cr
      -- 
    cp_elements(476) <= cp_elements(475);
    cr_10365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(476), ack => AND_u32_u32_2343_inst_req_1); -- 
    -- CP-element group 477 transition  output  bypass 
    -- predecessors 475 
    -- successors 478 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_tempx_x0x_xlcssax_xix_xi27_2340_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_tempx_x0x_xlcssax_xix_xi27_2340_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_tempx_x0x_xlcssax_xix_xi27_2340_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_tempx_x0x_xlcssax_xix_xi27_2340_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Sample/rr
      -- 
    cp_elements(477) <= cp_elements(475);
    rr_10360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => AND_u32_u32_2343_inst_req_0); -- 
    -- CP-element group 478 transition  input  bypass 
    -- predecessors 477 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Sample/ra
      -- 
    ra_10361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2343_inst_ack_0, ack => cp_elements(478)); -- 
    -- CP-element group 479 transition  input  bypass 
    -- predecessors 476 
    -- successors 487 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/AND_u32_u32_2343_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_112_2358_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_112_2358_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_112_2358_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_112_2358_update_completed_
      -- 
    ca_10366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2343_inst_ack_1, ack => cp_elements(479)); -- 
    -- CP-element group 480 transition  output  bypass 
    -- predecessors 475 
    -- successors 483 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Update/cr
      -- 
    cp_elements(480) <= cp_elements(475);
    cr_10383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(480), ack => SHL_u32_u32_2349_inst_req_1); -- 
    -- CP-element group 481 transition  output  bypass 
    -- predecessors 475 
    -- successors 482 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_expx_x0x_xlcssax_xix_xi26_2346_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_expx_x0x_xlcssax_xix_xi26_2346_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_expx_x0x_xlcssax_xix_xi26_2346_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_expx_x0x_xlcssax_xix_xi26_2346_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Sample/rr
      -- 
    cp_elements(481) <= cp_elements(475);
    rr_10378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(481), ack => SHL_u32_u32_2349_inst_req_0); -- 
    -- CP-element group 482 transition  input  bypass 
    -- predecessors 481 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Sample/ra
      -- 
    ra_10379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2349_inst_ack_0, ack => cp_elements(482)); -- 
    -- CP-element group 483 transition  input  output  bypass 
    -- predecessors 480 
    -- successors 485 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/SHL_u32_u32_2349_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_113_2352_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_113_2352_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_113_2352_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_113_2352_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Sample/rr
      -- 
    ca_10384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2349_inst_ack_1, ack => cp_elements(483)); -- 
    rr_10396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(483), ack => ADD_u32_u32_2355_inst_req_0); -- 
    -- CP-element group 484 transition  output  bypass 
    -- predecessors 475 
    -- successors 486 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Update/cr
      -- 
    cp_elements(484) <= cp_elements(475);
    cr_10401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => ADD_u32_u32_2355_inst_req_1); -- 
    -- CP-element group 485 transition  input  bypass 
    -- predecessors 483 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Sample/ra
      -- 
    ra_10397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2355_inst_ack_0, ack => cp_elements(485)); -- 
    -- CP-element group 486 transition  input  bypass 
    -- predecessors 484 
    -- successors 492 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/ADD_u32_u32_2355_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_114_2364_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_114_2364_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_114_2364_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_114_2364_update_completed_
      -- 
    ca_10402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2355_inst_ack_1, ack => cp_elements(486)); -- 
    -- CP-element group 487 join  transition  output  bypass 
    -- predecessors 479 489 
    -- successors 490 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Sample/rr
      -- 
    cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(479) & cp_elements(489);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(487), clk => clk, reset => reset); --
    end block;
    rr_10418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(487), ack => OR_u32_u32_2360_inst_req_0); -- 
    -- CP-element group 488 transition  output  bypass 
    -- predecessors 475 
    -- successors 491 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Update/cr
      -- 
    cp_elements(488) <= cp_elements(475);
    cr_10423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(488), ack => OR_u32_u32_2360_inst_req_1); -- 
    -- CP-element group 489 transition  bypass 
    -- predecessors 475 
    -- successors 487 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_63_2359_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_63_2359_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_63_2359_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_63_2359_update_completed_
      -- 
    cp_elements(489) <= cp_elements(475);
    -- CP-element group 490 transition  input  bypass 
    -- predecessors 487 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Sample/ra
      -- 
    ra_10419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2360_inst_ack_0, ack => cp_elements(490)); -- 
    -- CP-element group 491 transition  input  bypass 
    -- predecessors 488 
    -- successors 492 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2360_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_115_2363_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_115_2363_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_115_2363_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_115_2363_update_completed_
      -- 
    ca_10424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2360_inst_ack_1, ack => cp_elements(491)); -- 
    -- CP-element group 492 join  transition  output  bypass 
    -- predecessors 486 491 
    -- successors 494 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Sample/rr
      -- 
    cp_element_group_492: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_492"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(486) & cp_elements(491);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(492), clk => clk, reset => reset); --
    end block;
    rr_10440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(492), ack => OR_u32_u32_2365_inst_req_0); -- 
    -- CP-element group 493 transition  output  bypass 
    -- predecessors 475 
    -- successors 495 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Update/cr
      -- 
    cp_elements(493) <= cp_elements(475);
    cr_10445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(493), ack => OR_u32_u32_2365_inst_req_1); -- 
    -- CP-element group 494 transition  input  bypass 
    -- predecessors 492 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Sample/ra
      -- 
    ra_10441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2365_inst_ack_0, ack => cp_elements(494)); -- 
    -- CP-element group 495 transition  input  output  bypass 
    -- predecessors 493 
    -- successors 497 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_116_2368_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/OR_u32_u32_2365_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_116_2368_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_116_2368_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/R_iNsTr_116_2368_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Sample/rr
      -- 
    ca_10446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2365_inst_ack_1, ack => cp_elements(495)); -- 
    rr_10458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(495), ack => type_cast_2369_inst_req_0); -- 
    -- CP-element group 496 transition  output  bypass 
    -- predecessors 475 
    -- successors 498 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Update/cr
      -- 
    cp_elements(496) <= cp_elements(475);
    cr_10463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => type_cast_2369_inst_req_1); -- 
    -- CP-element group 497 transition  input  bypass 
    -- predecessors 495 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Sample/ra
      -- 
    ra_10459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2369_inst_ack_0, ack => cp_elements(497)); -- 
    -- CP-element group 498 fork  transition  place  input  bypass 
    -- predecessors 496 
    -- successors 1558 1560 
    -- members (11) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2344_to_assign_stmt_2370/type_cast_2369_Update/ca
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/$entry
      -- 
    ca_10464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2369_inst_ack_1, ack => cp_elements(498)); -- 
    -- CP-element group 499 fork  transition  bypass 
    -- predecessors 1565 
    -- successors 501 502 503 506 510 511 514 515 518 519 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/$entry
      -- 
    cp_elements(499) <= cp_elements(1565);
    -- CP-element group 500 join  transition  output  bypass 
    -- predecessors 502 503 
    -- successors 504 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Sample/rr
      -- 
    cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_500"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(502) & cp_elements(503);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(500), clk => clk, reset => reset); --
    end block;
    rr_10483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ADD_f32_f32_2384_inst_req_0); -- 
    -- CP-element group 501 transition  output  bypass 
    -- predecessors 499 
    -- successors 505 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Update/cr
      -- 
    cp_elements(501) <= cp_elements(499);
    cr_10488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => ADD_f32_f32_2384_inst_req_1); -- 
    -- CP-element group 502 transition  bypass 
    -- predecessors 499 
    -- successors 500 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_46_2382_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_46_2382_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_46_2382_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_46_2382_update_completed_
      -- 
    cp_elements(502) <= cp_elements(499);
    -- CP-element group 503 transition  bypass 
    -- predecessors 499 
    -- successors 500 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_10_2383_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_10_2383_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_10_2383_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_10_2383_update_completed_
      -- 
    cp_elements(503) <= cp_elements(499);
    -- CP-element group 504 transition  input  bypass 
    -- predecessors 500 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Sample/ra
      -- 
    ra_10484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2384_inst_ack_0, ack => cp_elements(504)); -- 
    -- CP-element group 505 transition  input  output  bypass 
    -- predecessors 501 
    -- successors 507 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2384_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_47_2387_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_47_2387_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_47_2387_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_47_2387_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Sample/rr
      -- 
    ca_10489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2384_inst_ack_1, ack => cp_elements(505)); -- 
    rr_10501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => MUL_f32_f32_2390_inst_req_0); -- 
    -- CP-element group 506 transition  output  bypass 
    -- predecessors 499 
    -- successors 508 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Update/cr
      -- 
    cp_elements(506) <= cp_elements(499);
    cr_10506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => MUL_f32_f32_2390_inst_req_1); -- 
    -- CP-element group 507 transition  input  bypass 
    -- predecessors 505 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Sample/ra
      -- 
    ra_10502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2390_inst_ack_0, ack => cp_elements(507)); -- 
    -- CP-element group 508 transition  input  bypass 
    -- predecessors 506 
    -- successors 509 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/MUL_f32_f32_2390_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_48_2393_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_48_2393_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_48_2393_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_iNsTr_48_2393_update_completed_
      -- 
    ca_10507_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2390_inst_ack_1, ack => cp_elements(508)); -- 
    -- CP-element group 509 join  transition  output  bypass 
    -- predecessors 508 511 
    -- successors 512 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Sample/rr
      -- 
    cp_element_group_509: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_509"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(508) & cp_elements(511);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(509), clk => clk, reset => reset); --
    end block;
    rr_10523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ADD_f32_f32_2395_inst_req_0); -- 
    -- CP-element group 510 transition  output  bypass 
    -- predecessors 499 
    -- successors 513 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Update/cr
      -- 
    cp_elements(510) <= cp_elements(499);
    cr_10528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(510), ack => ADD_f32_f32_2395_inst_req_1); -- 
    -- CP-element group 511 transition  bypass 
    -- predecessors 499 
    -- successors 509 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_theta_prevx_x0_2394_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_theta_prevx_x0_2394_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_theta_prevx_x0_2394_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_theta_prevx_x0_2394_update_completed_
      -- 
    cp_elements(511) <= cp_elements(499);
    -- CP-element group 512 transition  input  bypass 
    -- predecessors 509 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Sample/ra
      -- 
    ra_10524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2395_inst_ack_0, ack => cp_elements(512)); -- 
    -- CP-element group 513 transition  input  bypass 
    -- predecessors 510 
    -- successors 522 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/ADD_f32_f32_2395_Update/ca
      -- 
    ca_10529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2395_inst_ack_1, ack => cp_elements(513)); -- 
    -- CP-element group 514 transition  output  bypass 
    -- predecessors 499 
    -- successors 517 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Update/cr
      -- 
    cp_elements(514) <= cp_elements(499);
    cr_10546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => type_cast_2399_inst_req_1); -- 
    -- CP-element group 515 transition  output  bypass 
    -- predecessors 499 
    -- successors 516 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2398_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2398_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2398_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2398_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Sample/rr
      -- 
    cp_elements(515) <= cp_elements(499);
    rr_10541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => type_cast_2399_inst_req_0); -- 
    -- CP-element group 516 transition  input  bypass 
    -- predecessors 515 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Sample/ra
      -- 
    ra_10542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_0, ack => cp_elements(516)); -- 
    -- CP-element group 517 transition  input  bypass 
    -- predecessors 514 
    -- successors 522 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/type_cast_2399_Update/ca
      -- 
    ca_10547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_1, ack => cp_elements(517)); -- 
    -- CP-element group 518 transition  output  bypass 
    -- predecessors 499 
    -- successors 521 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Update/cr
      -- 
    cp_elements(518) <= cp_elements(499);
    cr_10564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(518), ack => EQ_f32_u1_2405_inst_req_1); -- 
    -- CP-element group 519 transition  output  bypass 
    -- predecessors 499 
    -- successors 520 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2402_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2402_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2402_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/R_torque_refx_x0_2402_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Sample/rr
      -- 
    cp_elements(519) <= cp_elements(499);
    rr_10559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => EQ_f32_u1_2405_inst_req_0); -- 
    -- CP-element group 520 transition  input  bypass 
    -- predecessors 519 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Sample/ra
      -- 
    ra_10560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2405_inst_ack_0, ack => cp_elements(520)); -- 
    -- CP-element group 521 transition  input  bypass 
    -- predecessors 518 
    -- successors 522 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/EQ_f32_u1_2405_Update/ca
      -- 
    ca_10565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2405_inst_ack_1, ack => cp_elements(521)); -- 
    -- CP-element group 522 join  transition  bypass 
    -- predecessors 513 517 521 
    -- successors 26 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406/$exit
      -- 
    cp_element_group_522: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_522"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(513) & cp_elements(517) & cp_elements(521);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(522), clk => clk, reset => reset); --
    end block;
    -- CP-element group 523 transition  place  dead  bypass 
    -- predecessors 26 
    -- successors 27 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2413__entry__
      -- 	branch_block_stmt_1659/if_stmt_2407__exit__
      -- 	branch_block_stmt_1659/if_stmt_2407_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2407_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2407_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2413_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2413_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2413_dead_link/dead_transition
      -- 
    cp_elements(523) <= false;
    -- CP-element group 524 transition  output  bypass 
    -- predecessors 26 
    -- successors 525 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2407_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2407_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2407_eval_test/branch_req
      -- 
    cp_elements(524) <= cp_elements(26);
    branch_req_10573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => if_stmt_2407_branch_req_0); -- 
    -- CP-element group 525 branch  place  bypass 
    -- predecessors 524 
    -- successors 526 528 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_50_2408_place
      -- 
    cp_elements(525) <= cp_elements(524);
    -- CP-element group 526 transition  bypass 
    -- predecessors 525 
    -- successors 527 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2407_if_link/$entry
      -- 
    cp_elements(526) <= cp_elements(525);
    -- CP-element group 527 fork  transition  place  input  bypass 
    -- predecessors 526 
    -- successors 1875 1876 
    -- members (8) 
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit
      -- 	branch_block_stmt_1659/if_stmt_2407_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2407_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/$entry
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/$entry
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/$entry
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/$entry
      -- 
    if_choice_transition_10578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2407_branch_ack_1, ack => cp_elements(527)); -- 
    -- CP-element group 528 transition  bypass 
    -- predecessors 525 
    -- successors 529 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2407_else_link/$entry
      -- 
    cp_elements(528) <= cp_elements(525);
    -- CP-element group 529 transition  place  input  bypass 
    -- predecessors 528 
    -- successors 27 
    -- members (9) 
      -- 	branch_block_stmt_1659/omega_calcx_xexit_bb_27
      -- 	branch_block_stmt_1659/if_stmt_2407_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2407_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/merge_stmt_2413_PhiReqMerge
      -- 	branch_block_stmt_1659/omega_calcx_xexit_bb_27_PhiReq/$entry
      -- 	branch_block_stmt_1659/omega_calcx_xexit_bb_27_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2413_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2413_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2413_PhiAck/dummy
      -- 
    else_choice_transition_10582_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2407_branch_ack_0, ack => cp_elements(529)); -- 
    -- CP-element group 530 fork  transition  bypass 
    -- predecessors 27 
    -- successors 531 532 535 538 539 542 545 546 549 552 555 556 559 562 566 567 568 571 575 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/$entry
      -- 
    cp_elements(530) <= cp_elements(27);
    -- CP-element group 531 transition  output  bypass 
    -- predecessors 530 
    -- successors 534 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Update/cr
      -- 
    cp_elements(531) <= cp_elements(530);
    cr_10604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(531), ack => LSHR_u32_u32_2418_inst_req_1); -- 
    -- CP-element group 532 transition  output  bypass 
    -- predecessors 530 
    -- successors 533 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2415_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2415_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2415_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2415_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Sample/rr
      -- 
    cp_elements(532) <= cp_elements(530);
    rr_10599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => LSHR_u32_u32_2418_inst_req_0); -- 
    -- CP-element group 533 transition  input  bypass 
    -- predecessors 532 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Sample/ra
      -- 
    ra_10600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2418_inst_ack_0, ack => cp_elements(533)); -- 
    -- CP-element group 534 transition  input  output  bypass 
    -- predecessors 531 
    -- successors 536 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2418_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_76_2421_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_76_2421_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_76_2421_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_76_2421_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Sample/rr
      -- 
    ca_10605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2418_inst_ack_1, ack => cp_elements(534)); -- 
    rr_10617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => AND_u32_u32_2424_inst_req_0); -- 
    -- CP-element group 535 transition  output  bypass 
    -- predecessors 530 
    -- successors 537 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Update/cr
      -- 
    cp_elements(535) <= cp_elements(530);
    cr_10622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => AND_u32_u32_2424_inst_req_1); -- 
    -- CP-element group 536 transition  input  bypass 
    -- predecessors 534 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Sample/ra
      -- 
    ra_10618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2424_inst_ack_0, ack => cp_elements(536)); -- 
    -- CP-element group 537 transition  input  bypass 
    -- predecessors 535 
    -- successors 574 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2424_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_77_2486_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_77_2486_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_77_2486_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_77_2486_update_completed_
      -- 
    ca_10623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2424_inst_ack_1, ack => cp_elements(537)); -- 
    -- CP-element group 538 transition  output  bypass 
    -- predecessors 530 
    -- successors 541 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Update/cr
      -- 
    cp_elements(538) <= cp_elements(530);
    cr_10640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => LSHR_u32_u32_2430_inst_req_1); -- 
    -- CP-element group 539 transition  output  bypass 
    -- predecessors 530 
    -- successors 540 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2427_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2427_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2427_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2427_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Sample/rr
      -- 
    cp_elements(539) <= cp_elements(530);
    rr_10635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(539), ack => LSHR_u32_u32_2430_inst_req_0); -- 
    -- CP-element group 540 transition  input  bypass 
    -- predecessors 539 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Sample/ra
      -- 
    ra_10636_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2430_inst_ack_0, ack => cp_elements(540)); -- 
    -- CP-element group 541 transition  input  output  bypass 
    -- predecessors 538 
    -- successors 543 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2430_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_78_2433_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_78_2433_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_78_2433_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_78_2433_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Sample/rr
      -- 
    ca_10641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2430_inst_ack_1, ack => cp_elements(541)); -- 
    rr_10653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => AND_u32_u32_2436_inst_req_0); -- 
    -- CP-element group 542 transition  output  bypass 
    -- predecessors 530 
    -- successors 544 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Update/cr
      -- 
    cp_elements(542) <= cp_elements(530);
    cr_10658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(542), ack => AND_u32_u32_2436_inst_req_1); -- 
    -- CP-element group 543 transition  input  bypass 
    -- predecessors 541 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Sample/ra
      -- 
    ra_10654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2436_inst_ack_0, ack => cp_elements(543)); -- 
    -- CP-element group 544 transition  input  bypass 
    -- predecessors 542 
    -- successors 574 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2436_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_79_2487_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_79_2487_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_79_2487_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_79_2487_update_completed_
      -- 
    ca_10659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2436_inst_ack_1, ack => cp_elements(544)); -- 
    -- CP-element group 545 transition  output  bypass 
    -- predecessors 530 
    -- successors 548 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Update/cr
      -- 
    cp_elements(545) <= cp_elements(530);
    cr_10676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => SHL_u32_u32_2442_inst_req_1); -- 
    -- CP-element group 546 transition  output  bypass 
    -- predecessors 530 
    -- successors 547 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2439_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2439_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2439_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2439_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Sample/rr
      -- 
    cp_elements(546) <= cp_elements(530);
    rr_10671_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(546), ack => SHL_u32_u32_2442_inst_req_0); -- 
    -- CP-element group 547 transition  input  bypass 
    -- predecessors 546 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Sample/ra
      -- 
    ra_10672_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2442_inst_ack_0, ack => cp_elements(547)); -- 
    -- CP-element group 548 transition  input  output  bypass 
    -- predecessors 545 
    -- successors 550 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SHL_u32_u32_2442_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_80_2445_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_80_2445_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_80_2445_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_80_2445_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Sample/rr
      -- 
    ca_10677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2442_inst_ack_1, ack => cp_elements(548)); -- 
    rr_10689_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => AND_u32_u32_2448_inst_req_0); -- 
    -- CP-element group 549 transition  output  bypass 
    -- predecessors 530 
    -- successors 551 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Update/cr
      -- 
    cp_elements(549) <= cp_elements(530);
    cr_10694_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => AND_u32_u32_2448_inst_req_1); -- 
    -- CP-element group 550 transition  input  bypass 
    -- predecessors 548 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Sample/ra
      -- 
    ra_10690_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2448_inst_ack_0, ack => cp_elements(550)); -- 
    -- CP-element group 551 transition  input  output  bypass 
    -- predecessors 549 
    -- successors 553 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2448_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_81_2451_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_81_2451_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_81_2451_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_81_2451_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Sample/rr
      -- 
    ca_10695_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2448_inst_ack_1, ack => cp_elements(551)); -- 
    rr_10707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(551), ack => OR_u32_u32_2454_inst_req_0); -- 
    -- CP-element group 552 transition  output  bypass 
    -- predecessors 530 
    -- successors 554 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Update/cr
      -- 
    cp_elements(552) <= cp_elements(530);
    cr_10712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => OR_u32_u32_2454_inst_req_1); -- 
    -- CP-element group 553 transition  input  bypass 
    -- predecessors 551 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Sample/ra
      -- 
    ra_10708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2454_inst_ack_0, ack => cp_elements(553)); -- 
    -- CP-element group 554 transition  input  bypass 
    -- predecessors 552 
    -- successors 578 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2454_Update/ca
      -- 
    ca_10713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2454_inst_ack_1, ack => cp_elements(554)); -- 
    -- CP-element group 555 transition  output  bypass 
    -- predecessors 530 
    -- successors 558 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Update/cr
      -- 
    cp_elements(555) <= cp_elements(530);
    cr_10730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(555), ack => LSHR_u32_u32_2460_inst_req_1); -- 
    -- CP-element group 556 transition  output  bypass 
    -- predecessors 530 
    -- successors 557 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2457_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2457_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2457_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2457_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Sample/rr
      -- 
    cp_elements(556) <= cp_elements(530);
    rr_10725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => LSHR_u32_u32_2460_inst_req_0); -- 
    -- CP-element group 557 transition  input  bypass 
    -- predecessors 556 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Sample/ra
      -- 
    ra_10726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2460_inst_ack_0, ack => cp_elements(557)); -- 
    -- CP-element group 558 transition  input  output  bypass 
    -- predecessors 555 
    -- successors 560 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/LSHR_u32_u32_2460_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_83_2463_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_83_2463_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_83_2463_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_83_2463_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Sample/rr
      -- 
    ca_10731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2460_inst_ack_1, ack => cp_elements(558)); -- 
    rr_10743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(558), ack => AND_u32_u32_2466_inst_req_0); -- 
    -- CP-element group 559 transition  output  bypass 
    -- predecessors 530 
    -- successors 561 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Update/cr
      -- 
    cp_elements(559) <= cp_elements(530);
    cr_10748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => AND_u32_u32_2466_inst_req_1); -- 
    -- CP-element group 560 transition  input  bypass 
    -- predecessors 558 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Sample/ra
      -- 
    ra_10744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2466_inst_ack_0, ack => cp_elements(560)); -- 
    -- CP-element group 561 transition  input  output  bypass 
    -- predecessors 559 
    -- successors 563 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2466_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_84_2469_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_84_2469_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_84_2469_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_84_2469_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Sample/rr
      -- 
    ca_10749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2466_inst_ack_1, ack => cp_elements(561)); -- 
    rr_10761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => OR_u32_u32_2472_inst_req_0); -- 
    -- CP-element group 562 transition  output  bypass 
    -- predecessors 530 
    -- successors 564 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Update/cr
      -- 
    cp_elements(562) <= cp_elements(530);
    cr_10766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(562), ack => OR_u32_u32_2472_inst_req_1); -- 
    -- CP-element group 563 transition  input  bypass 
    -- predecessors 561 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Sample/ra
      -- 
    ra_10762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2472_inst_ack_0, ack => cp_elements(563)); -- 
    -- CP-element group 564 transition  input  bypass 
    -- predecessors 562 
    -- successors 578 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/OR_u32_u32_2472_Update/ca
      -- 
    ca_10767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2472_inst_ack_1, ack => cp_elements(564)); -- 
    -- CP-element group 565 join  transition  output  bypass 
    -- predecessors 567 568 
    -- successors 569 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Sample/rr
      -- 
    cp_element_group_565: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_565"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(567) & cp_elements(568);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(565), clk => clk, reset => reset); --
    end block;
    rr_10783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => XOR_u32_u32_2477_inst_req_0); -- 
    -- CP-element group 566 transition  output  bypass 
    -- predecessors 530 
    -- successors 570 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Update/cr
      -- 
    cp_elements(566) <= cp_elements(530);
    cr_10788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => XOR_u32_u32_2477_inst_req_1); -- 
    -- CP-element group 567 transition  bypass 
    -- predecessors 530 
    -- successors 565 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2475_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2475_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2475_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp10x_xix_xi_2475_update_completed_
      -- 
    cp_elements(567) <= cp_elements(530);
    -- CP-element group 568 transition  bypass 
    -- predecessors 530 
    -- successors 565 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2476_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2476_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2476_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_tmp6x_xix_xi2_2476_update_completed_
      -- 
    cp_elements(568) <= cp_elements(530);
    -- CP-element group 569 transition  input  bypass 
    -- predecessors 565 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Sample/ra
      -- 
    ra_10784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2477_inst_ack_0, ack => cp_elements(569)); -- 
    -- CP-element group 570 transition  input  output  bypass 
    -- predecessors 566 
    -- successors 572 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/XOR_u32_u32_2477_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_86_2480_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_86_2480_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_86_2480_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/R_iNsTr_86_2480_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Sample/rr
      -- 
    ca_10789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2477_inst_ack_1, ack => cp_elements(570)); -- 
    rr_10801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(570), ack => AND_u32_u32_2483_inst_req_0); -- 
    -- CP-element group 571 transition  output  bypass 
    -- predecessors 530 
    -- successors 573 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Update/cr
      -- 
    cp_elements(571) <= cp_elements(530);
    cr_10806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => AND_u32_u32_2483_inst_req_1); -- 
    -- CP-element group 572 transition  input  bypass 
    -- predecessors 570 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Sample/ra
      -- 
    ra_10802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2483_inst_ack_0, ack => cp_elements(572)); -- 
    -- CP-element group 573 transition  input  bypass 
    -- predecessors 571 
    -- successors 578 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/AND_u32_u32_2483_Update/ca
      -- 
    ca_10807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2483_inst_ack_1, ack => cp_elements(573)); -- 
    -- CP-element group 574 join  transition  output  bypass 
    -- predecessors 537 544 
    -- successors 576 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Sample/rr
      -- 
    cp_element_group_574: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_574"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(537) & cp_elements(544);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(574), clk => clk, reset => reset); --
    end block;
    rr_10823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => SUB_u32_u32_2488_inst_req_0); -- 
    -- CP-element group 575 transition  output  bypass 
    -- predecessors 530 
    -- successors 577 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Update/cr
      -- 
    cp_elements(575) <= cp_elements(530);
    cr_10828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => SUB_u32_u32_2488_inst_req_1); -- 
    -- CP-element group 576 transition  input  bypass 
    -- predecessors 574 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Sample/ra
      -- 
    ra_10824_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2488_inst_ack_0, ack => cp_elements(576)); -- 
    -- CP-element group 577 transition  input  bypass 
    -- predecessors 575 
    -- successors 578 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/SUB_u32_u32_2488_Update/ca
      -- 
    ca_10829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2488_inst_ack_1, ack => cp_elements(577)); -- 
    -- CP-element group 578 join  transition  bypass 
    -- predecessors 554 564 573 577 
    -- successors 28 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2419_to_assign_stmt_2489/$exit
      -- 
    cp_element_group_578: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_578"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= cp_elements(554) & cp_elements(564) & cp_elements(573) & cp_elements(577);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(578), clk => clk, reset => reset); --
    end block;
    -- CP-element group 579 transition  place  dead  bypass 
    -- predecessors 28 
    -- successors 29 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2500__entry__
      -- 	branch_block_stmt_1659/switch_stmt_2490__exit__
      -- 	branch_block_stmt_1659/switch_stmt_2490_dead_link/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490_dead_link/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2500_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2500_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2500_dead_link/dead_transition
      -- 
    cp_elements(579) <= false;
    -- CP-element group 580 place  bypass 
    -- predecessors 28 
    -- successors 581 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check_place__
      -- 
    cp_elements(580) <= cp_elements(28);
    -- CP-element group 581 fork  transition  bypass 
    -- predecessors 580 
    -- successors 582 588 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/$entry
      -- 
    cp_elements(581) <= cp_elements(580);
    -- CP-element group 582 fork  transition  bypass 
    -- predecessors 581 
    -- successors 583 585 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/$entry
      -- 
    cp_elements(582) <= cp_elements(581);
    -- CP-element group 583 transition  output  bypass 
    -- predecessors 582 
    -- successors 584 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Sample/rr
      -- 
    cp_elements(583) <= cp_elements(582);
    rr_10847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(583), ack => switch_stmt_2490_select_expr_0_req_0); -- 
    -- CP-element group 584 transition  input  bypass 
    -- predecessors 583 
    -- successors 587 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Sample/ra
      -- 
    ra_10848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_select_expr_0_ack_0, ack => cp_elements(584)); -- 
    -- CP-element group 585 transition  output  bypass 
    -- predecessors 582 
    -- successors 586 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Update/cr
      -- 
    cp_elements(585) <= cp_elements(582);
    cr_10852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(585), ack => switch_stmt_2490_select_expr_0_req_1); -- 
    -- CP-element group 586 transition  input  bypass 
    -- predecessors 585 
    -- successors 587 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/Update/ca
      -- 
    ca_10853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_select_expr_0_ack_1, ack => cp_elements(586)); -- 
    -- CP-element group 587 join  transition  output  bypass 
    -- predecessors 584 586 
    -- successors 594 
    -- members (3) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_0/cmp
      -- 
    cp_element_group_587: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_587"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(584) & cp_elements(586);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(587), clk => clk, reset => reset); --
    end block;
    cmp_10854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => switch_stmt_2490_branch_0_req_0); -- 
    -- CP-element group 588 fork  transition  bypass 
    -- predecessors 581 
    -- successors 589 591 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/$entry
      -- 
    cp_elements(588) <= cp_elements(581);
    -- CP-element group 589 transition  output  bypass 
    -- predecessors 588 
    -- successors 590 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Sample/rr
      -- 
    cp_elements(589) <= cp_elements(588);
    rr_10864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(589), ack => switch_stmt_2490_select_expr_1_req_0); -- 
    -- CP-element group 590 transition  input  bypass 
    -- predecessors 589 
    -- successors 593 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Sample/ra
      -- 
    ra_10865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_select_expr_1_ack_0, ack => cp_elements(590)); -- 
    -- CP-element group 591 transition  output  bypass 
    -- predecessors 588 
    -- successors 592 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Update/cr
      -- 
    cp_elements(591) <= cp_elements(588);
    cr_10869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => switch_stmt_2490_select_expr_1_req_1); -- 
    -- CP-element group 592 transition  input  bypass 
    -- predecessors 591 
    -- successors 593 
    -- members (2) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/Update/ca
      -- 
    ca_10870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_select_expr_1_ack_1, ack => cp_elements(592)); -- 
    -- CP-element group 593 join  transition  output  bypass 
    -- predecessors 590 592 
    -- successors 594 
    -- members (3) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/condition_1/cmp
      -- 
    cp_element_group_593: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_593"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(590) & cp_elements(592);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(593), clk => clk, reset => reset); --
    end block;
    cmp_10871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => switch_stmt_2490_branch_1_req_0); -- 
    -- CP-element group 594 join  transition  output  bypass 
    -- predecessors 587 593 
    -- successors 595 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__condition_check__/$exit
      -- 
    cp_element_group_594: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_594"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(587) & cp_elements(593);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(594), clk => clk, reset => reset); --
    end block;
    Xexit_10837_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(594), ack => switch_stmt_2490_branch_default_req_0); -- 
    -- CP-element group 595 branch  place  bypass 
    -- predecessors 594 
    -- successors 596 598 600 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490__select__
      -- 
    cp_elements(595) <= cp_elements(594);
    -- CP-element group 596 transition  bypass 
    -- predecessors 595 
    -- successors 597 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_0/$entry
      -- 
    cp_elements(596) <= cp_elements(595);
    -- CP-element group 597 fork  transition  place  input  bypass 
    -- predecessors 596 
    -- successors 1720 1721 
    -- members (8) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_0/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_0/ack1
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/$entry
      -- 
    ack1_10876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_branch_0_ack_1, ack => cp_elements(597)); -- 
    -- CP-element group 598 transition  bypass 
    -- predecessors 595 
    -- successors 599 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_1/$entry
      -- 
    cp_elements(598) <= cp_elements(595);
    -- CP-element group 599 fork  transition  place  input  bypass 
    -- predecessors 598 
    -- successors 1731 1735 
    -- members (6) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_1/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_1/ack1
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/$entry
      -- 
    ack1_10881_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_branch_1_ack_1, ack => cp_elements(599)); -- 
    -- CP-element group 600 transition  bypass 
    -- predecessors 595 
    -- successors 601 
    -- members (1) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_default/$entry
      -- 
    cp_elements(600) <= cp_elements(595);
    -- CP-element group 601 transition  place  input  bypass 
    -- predecessors 600 
    -- successors 29 
    -- members (9) 
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_default/$exit
      -- 	branch_block_stmt_1659/switch_stmt_2490_choice_default/ack0
      -- 	branch_block_stmt_1659/bb_27_bbx_xnph7x_xix_xix_xix_xpreheader
      -- 	branch_block_stmt_1659/merge_stmt_2500_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_27_bbx_xnph7x_xix_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_27_bbx_xnph7x_xix_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2500_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2500_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2500_PhiAck/dummy
      -- 
    ack0_10886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_2490_branch_default_ack_0, ack => cp_elements(601)); -- 
    -- CP-element group 602 fork  transition  bypass 
    -- predecessors 30 
    -- successors 603 604 608 609 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/$entry
      -- 
    cp_elements(602) <= cp_elements(30);
    -- CP-element group 603 transition  output  bypass 
    -- predecessors 602 
    -- successors 606 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Update/cr
      -- 
    cp_elements(603) <= cp_elements(602);
    cr_10907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(603), ack => LSHR_u32_u32_2521_inst_req_1); -- 
    -- CP-element group 604 transition  output  bypass 
    -- predecessors 602 
    -- successors 605 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_xx_x016x_xix_xix_xi_2518_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_xx_x016x_xix_xix_xi_2518_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_xx_x016x_xix_xix_xi_2518_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_xx_x016x_xix_xix_xi_2518_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Sample/rr
      -- 
    cp_elements(604) <= cp_elements(602);
    rr_10902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => LSHR_u32_u32_2521_inst_req_0); -- 
    -- CP-element group 605 transition  input  bypass 
    -- predecessors 604 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Sample/ra
      -- 
    ra_10903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2521_inst_ack_0, ack => cp_elements(605)); -- 
    -- CP-element group 606 transition  input  bypass 
    -- predecessors 603 
    -- successors 607 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/LSHR_u32_u32_2521_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_125_2524_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_125_2524_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_125_2524_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_125_2524_update_completed_
      -- 
    ca_10908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_2521_inst_ack_1, ack => cp_elements(606)); -- 
    -- CP-element group 607 join  transition  output  bypass 
    -- predecessors 606 609 
    -- successors 610 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Sample/rr
      -- 
    cp_element_group_607: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_607"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(606) & cp_elements(609);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(607), clk => clk, reset => reset); --
    end block;
    rr_10924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(607), ack => UGT_u32_u1_2526_inst_req_0); -- 
    -- CP-element group 608 transition  output  bypass 
    -- predecessors 602 
    -- successors 611 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Update/cr
      -- 
    cp_elements(608) <= cp_elements(602);
    cr_10929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(608), ack => UGT_u32_u1_2526_inst_req_1); -- 
    -- CP-element group 609 transition  bypass 
    -- predecessors 602 
    -- successors 607 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_85_2525_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_85_2525_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_85_2525_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/R_iNsTr_85_2525_update_completed_
      -- 
    cp_elements(609) <= cp_elements(602);
    -- CP-element group 610 transition  input  bypass 
    -- predecessors 607 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Sample/ra
      -- 
    ra_10925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2526_inst_ack_0, ack => cp_elements(610)); -- 
    -- CP-element group 611 branch  transition  place  input  bypass 
    -- predecessors 608 
    -- successors 612 613 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527__exit__
      -- 	branch_block_stmt_1659/if_stmt_2528__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2522_to_assign_stmt_2527/UGT_u32_u1_2526_Update/ca
      -- 
    ca_10930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_2526_inst_ack_1, ack => cp_elements(611)); -- 
    -- CP-element group 612 transition  place  dead  bypass 
    -- predecessors 611 
    -- successors 31 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2534__entry__
      -- 	branch_block_stmt_1659/if_stmt_2528__exit__
      -- 	branch_block_stmt_1659/if_stmt_2528_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2528_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2528_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2534_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2534_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2534_dead_link/dead_transition
      -- 
    cp_elements(612) <= false;
    -- CP-element group 613 transition  output  bypass 
    -- predecessors 611 
    -- successors 614 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2528_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2528_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2528_eval_test/branch_req
      -- 
    cp_elements(613) <= cp_elements(611);
    branch_req_10938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => if_stmt_2528_branch_req_0); -- 
    -- CP-element group 614 branch  place  bypass 
    -- predecessors 613 
    -- successors 615 617 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_126_2529_place
      -- 
    cp_elements(614) <= cp_elements(613);
    -- CP-element group 615 transition  bypass 
    -- predecessors 614 
    -- successors 616 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2528_if_link/$entry
      -- 
    cp_elements(615) <= cp_elements(614);
    -- CP-element group 616 transition  place  input  bypass 
    -- predecessors 615 
    -- successors 31 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2528_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2528_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader
      -- 	branch_block_stmt_1659/merge_stmt_2534_PhiReqMerge
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_bbx_xnphx_xix_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2534_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2534_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2534_PhiAck/dummy
      -- 
    if_choice_transition_10943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2528_branch_ack_1, ack => cp_elements(616)); -- 
    -- CP-element group 617 transition  bypass 
    -- predecessors 614 
    -- successors 618 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2528_else_link/$entry
      -- 
    cp_elements(617) <= cp_elements(614);
    -- CP-element group 618 transition  place  input  bypass 
    -- predecessors 617 
    -- successors 1671 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2528_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2528_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi
      -- 
    else_choice_transition_10947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2528_branch_ack_0, ack => cp_elements(618)); -- 
    -- CP-element group 619 fork  transition  bypass 
    -- predecessors 32 
    -- successors 620 621 624 625 629 630 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/$entry
      -- 
    cp_elements(619) <= cp_elements(32);
    -- CP-element group 620 transition  output  bypass 
    -- predecessors 619 
    -- successors 623 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Update/cr
      -- 
    cp_elements(620) <= cp_elements(619);
    cr_10969_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(620), ack => SHL_u32_u32_2555_inst_req_1); -- 
    -- CP-element group 621 transition  output  bypass 
    -- predecessors 619 
    -- successors 622 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_shifted_divisorx_x03x_xix_xix_xi_2552_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_shifted_divisorx_x03x_xix_xix_xi_2552_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_shifted_divisorx_x03x_xix_xix_xi_2552_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_shifted_divisorx_x03x_xix_xix_xi_2552_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Sample/rr
      -- 
    cp_elements(621) <= cp_elements(619);
    rr_10964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => SHL_u32_u32_2555_inst_req_0); -- 
    -- CP-element group 622 transition  input  bypass 
    -- predecessors 621 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Sample/ra
      -- 
    ra_10965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2555_inst_ack_0, ack => cp_elements(622)); -- 
    -- CP-element group 623 transition  input  bypass 
    -- predecessors 620 
    -- successors 628 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2555_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_183_2564_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_183_2564_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_183_2564_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_183_2564_update_completed_
      -- 
    ca_10970_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2555_inst_ack_1, ack => cp_elements(623)); -- 
    -- CP-element group 624 transition  output  bypass 
    -- predecessors 619 
    -- successors 627 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Update/cr
      -- 
    cp_elements(624) <= cp_elements(619);
    cr_10987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(624), ack => SHL_u32_u32_2561_inst_req_1); -- 
    -- CP-element group 625 transition  output  bypass 
    -- predecessors 619 
    -- successors 626 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_curr_quotientx_x02x_xix_xix_xi_2558_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_curr_quotientx_x02x_xix_xix_xi_2558_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_curr_quotientx_x02x_xix_xix_xi_2558_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_curr_quotientx_x02x_xix_xix_xi_2558_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Sample/rr
      -- 
    cp_elements(625) <= cp_elements(619);
    rr_10982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(625), ack => SHL_u32_u32_2561_inst_req_0); -- 
    -- CP-element group 626 transition  input  bypass 
    -- predecessors 625 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Sample/ra
      -- 
    ra_10983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2561_inst_ack_0, ack => cp_elements(626)); -- 
    -- CP-element group 627 transition  input  bypass 
    -- predecessors 624 
    -- successors 633 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/SHL_u32_u32_2561_Update/ca
      -- 
    ca_10988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2561_inst_ack_1, ack => cp_elements(627)); -- 
    -- CP-element group 628 join  transition  output  bypass 
    -- predecessors 623 630 
    -- successors 631 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Sample/rr
      -- 
    cp_element_group_628: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_628"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(623) & cp_elements(630);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(628), clk => clk, reset => reset); --
    end block;
    rr_11004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(628), ack => ULT_u32_u1_2566_inst_req_0); -- 
    -- CP-element group 629 transition  output  bypass 
    -- predecessors 619 
    -- successors 632 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Update/cr
      -- 
    cp_elements(629) <= cp_elements(619);
    cr_11009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(629), ack => ULT_u32_u1_2566_inst_req_1); -- 
    -- CP-element group 630 transition  bypass 
    -- predecessors 619 
    -- successors 628 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_125_2565_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_125_2565_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_125_2565_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/R_iNsTr_125_2565_update_completed_
      -- 
    cp_elements(630) <= cp_elements(619);
    -- CP-element group 631 transition  input  bypass 
    -- predecessors 628 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Sample/ra
      -- 
    ra_11005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2566_inst_ack_0, ack => cp_elements(631)); -- 
    -- CP-element group 632 transition  input  bypass 
    -- predecessors 629 
    -- successors 633 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/ULT_u32_u1_2566_Update/ca
      -- 
    ca_11010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2566_inst_ack_1, ack => cp_elements(632)); -- 
    -- CP-element group 633 join  transition  bypass 
    -- predecessors 627 632 
    -- successors 33 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2556_to_assign_stmt_2567/$exit
      -- 
    cp_element_group_633: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_633"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(627) & cp_elements(632);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(633), clk => clk, reset => reset); --
    end block;
    -- CP-element group 634 transition  place  dead  bypass 
    -- predecessors 33 
    -- successors 34 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2568__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2574__entry__
      -- 	branch_block_stmt_1659/if_stmt_2568_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2568_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2568_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2574_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2574_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2574_dead_link/dead_transition
      -- 
    cp_elements(634) <= false;
    -- CP-element group 635 transition  output  bypass 
    -- predecessors 33 
    -- successors 636 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2568_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2568_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2568_eval_test/branch_req
      -- 
    cp_elements(635) <= cp_elements(33);
    branch_req_11018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(635), ack => if_stmt_2568_branch_req_0); -- 
    -- CP-element group 636 branch  place  bypass 
    -- predecessors 635 
    -- successors 637 639 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_185_2569_place
      -- 
    cp_elements(636) <= cp_elements(635);
    -- CP-element group 637 transition  bypass 
    -- predecessors 636 
    -- successors 638 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2568_if_link/$entry
      -- 
    cp_elements(637) <= cp_elements(636);
    -- CP-element group 638 transition  place  input  bypass 
    -- predecessors 637 
    -- successors 1609 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2568_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2568_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi
      -- 
    if_choice_transition_11023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2568_branch_ack_1, ack => cp_elements(638)); -- 
    -- CP-element group 639 transition  bypass 
    -- predecessors 636 
    -- successors 640 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2568_else_link/$entry
      -- 
    cp_elements(639) <= cp_elements(636);
    -- CP-element group 640 transition  place  input  bypass 
    -- predecessors 639 
    -- successors 1652 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2568_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2568_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit
      -- 
    else_choice_transition_11027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2568_branch_ack_0, ack => cp_elements(640)); -- 
    -- CP-element group 641 fork  transition  bypass 
    -- predecessors 35 
    -- successors 643 644 645 649 650 651 655 656 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/$entry
      -- 
    cp_elements(641) <= cp_elements(35);
    -- CP-element group 642 join  transition  output  bypass 
    -- predecessors 644 645 
    -- successors 646 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Sample/rr
      -- 
    cp_element_group_642: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_642"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(644) & cp_elements(645);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(642), clk => clk, reset => reset); --
    end block;
    rr_11048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => ADD_u32_u32_2603_inst_req_0); -- 
    -- CP-element group 643 transition  output  bypass 
    -- predecessors 641 
    -- successors 647 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Update/cr
      -- 
    cp_elements(643) <= cp_elements(641);
    cr_11053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => ADD_u32_u32_2603_inst_req_1); -- 
    -- CP-element group 644 transition  bypass 
    -- predecessors 641 
    -- successors 642 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_2601_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_2601_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_2601_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_curr_quotientx_x0x_xlcssax_xix_xix_xi_2601_update_completed_
      -- 
    cp_elements(644) <= cp_elements(641);
    -- CP-element group 645 transition  bypass 
    -- predecessors 641 
    -- successors 642 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_quotientx_x05x_xix_xix_xi_2602_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_quotientx_x05x_xix_xix_xi_2602_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_quotientx_x05x_xix_xix_xi_2602_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_quotientx_x05x_xix_xix_xi_2602_update_completed_
      -- 
    cp_elements(645) <= cp_elements(641);
    -- CP-element group 646 transition  input  bypass 
    -- predecessors 642 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Sample/ra
      -- 
    ra_11049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2603_inst_ack_0, ack => cp_elements(646)); -- 
    -- CP-element group 647 transition  input  bypass 
    -- predecessors 643 
    -- successors 659 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ADD_u32_u32_2603_Update/ca
      -- 
    ca_11054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2603_inst_ack_1, ack => cp_elements(647)); -- 
    -- CP-element group 648 join  transition  output  bypass 
    -- predecessors 650 651 
    -- successors 652 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Sample/rr
      -- 
    cp_element_group_648: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_648"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(650) & cp_elements(651);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(648), clk => clk, reset => reset); --
    end block;
    rr_11070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(648), ack => SUB_u32_u32_2608_inst_req_0); -- 
    -- CP-element group 649 transition  output  bypass 
    -- predecessors 641 
    -- successors 653 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Update/cr
      -- 
    cp_elements(649) <= cp_elements(641);
    cr_11075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(649), ack => SUB_u32_u32_2608_inst_req_1); -- 
    -- CP-element group 650 transition  bypass 
    -- predecessors 641 
    -- successors 648 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_xx_x016x_xix_xix_xi_2606_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_xx_x016x_xix_xix_xi_2606_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_xx_x016x_xix_xix_xi_2606_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_xx_x016x_xix_xix_xi_2606_update_completed_
      -- 
    cp_elements(650) <= cp_elements(641);
    -- CP-element group 651 transition  bypass 
    -- predecessors 641 
    -- successors 648 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_2607_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_2607_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_2607_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_shifted_divisorx_x0x_xlcssax_xix_xix_xi_2607_update_completed_
      -- 
    cp_elements(651) <= cp_elements(641);
    -- CP-element group 652 transition  input  bypass 
    -- predecessors 648 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Sample/ra
      -- 
    ra_11071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2608_inst_ack_0, ack => cp_elements(652)); -- 
    -- CP-element group 653 transition  input  bypass 
    -- predecessors 649 
    -- successors 654 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/SUB_u32_u32_2608_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_153_2611_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_153_2611_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_153_2611_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_153_2611_update_completed_
      -- 
    ca_11076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2608_inst_ack_1, ack => cp_elements(653)); -- 
    -- CP-element group 654 join  transition  output  bypass 
    -- predecessors 653 656 
    -- successors 657 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Sample/rr
      -- 
    cp_element_group_654: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_654"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(653) & cp_elements(656);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(654), clk => clk, reset => reset); --
    end block;
    rr_11092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ULT_u32_u1_2613_inst_req_0); -- 
    -- CP-element group 655 transition  output  bypass 
    -- predecessors 641 
    -- successors 658 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Update/cr
      -- 
    cp_elements(655) <= cp_elements(641);
    cr_11097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => ULT_u32_u1_2613_inst_req_1); -- 
    -- CP-element group 656 transition  bypass 
    -- predecessors 641 
    -- successors 654 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_85_2612_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_85_2612_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_85_2612_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/R_iNsTr_85_2612_update_completed_
      -- 
    cp_elements(656) <= cp_elements(641);
    -- CP-element group 657 transition  input  bypass 
    -- predecessors 654 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Sample/ra
      -- 
    ra_11093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2613_inst_ack_0, ack => cp_elements(657)); -- 
    -- CP-element group 658 transition  input  bypass 
    -- predecessors 655 
    -- successors 659 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/ULT_u32_u1_2613_Update/ca
      -- 
    ca_11098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_2613_inst_ack_1, ack => cp_elements(658)); -- 
    -- CP-element group 659 join  transition  bypass 
    -- predecessors 647 658 
    -- successors 36 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2604_to_assign_stmt_2614/$exit
      -- 
    cp_element_group_659: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_659"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(647) & cp_elements(658);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(659), clk => clk, reset => reset); --
    end block;
    -- CP-element group 660 transition  place  dead  bypass 
    -- predecessors 36 
    -- successors 37 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2615__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2621__entry__
      -- 	branch_block_stmt_1659/if_stmt_2615_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2615_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2615_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2621_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2621_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2621_dead_link/dead_transition
      -- 
    cp_elements(660) <= false;
    -- CP-element group 661 transition  output  bypass 
    -- predecessors 36 
    -- successors 662 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2615_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2615_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2615_eval_test/branch_req
      -- 
    cp_elements(661) <= cp_elements(36);
    branch_req_11106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(661), ack => if_stmt_2615_branch_req_0); -- 
    -- CP-element group 662 branch  place  bypass 
    -- predecessors 661 
    -- successors 663 665 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_154_2616_place
      -- 
    cp_elements(662) <= cp_elements(661);
    -- CP-element group 663 transition  bypass 
    -- predecessors 662 
    -- successors 664 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2615_if_link/$entry
      -- 
    cp_elements(663) <= cp_elements(662);
    -- CP-element group 664 fork  transition  place  input  bypass 
    -- predecessors 663 
    -- successors 1714 1716 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2615_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2615_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/$entry
      -- 
    if_choice_transition_11111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2615_branch_ack_1, ack => cp_elements(664)); -- 
    -- CP-element group 665 transition  bypass 
    -- predecessors 662 
    -- successors 666 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2615_else_link/$entry
      -- 
    cp_elements(665) <= cp_elements(662);
    -- CP-element group 666 transition  place  input  bypass 
    -- predecessors 665 
    -- successors 1584 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2615_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2615_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi
      -- 
    else_choice_transition_11115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2615_branch_ack_0, ack => cp_elements(666)); -- 
    -- CP-element group 667 fork  transition  bypass 
    -- predecessors 1755 
    -- successors 668 669 672 675 676 682 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/$entry
      -- 
    cp_elements(667) <= cp_elements(1755);
    -- CP-element group 668 transition  output  bypass 
    -- predecessors 667 
    -- successors 671 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_update_start_
      -- 
    cp_elements(668) <= cp_elements(667);
    cr_11137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => AND_u32_u32_2650_inst_req_1); -- 
    -- CP-element group 669 transition  output  bypass 
    -- predecessors 667 
    -- successors 670 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2647_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2647_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2647_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2647_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_sample_start_
      -- 
    cp_elements(669) <= cp_elements(667);
    rr_11132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(669), ack => AND_u32_u32_2650_inst_req_0); -- 
    -- CP-element group 670 transition  input  bypass 
    -- predecessors 669 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_sample_completed_
      -- 
    ra_11133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2650_inst_ack_0, ack => cp_elements(670)); -- 
    -- CP-element group 671 transition  input  output  bypass 
    -- predecessors 668 
    -- successors 673 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_104_2653_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_104_2653_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_104_2653_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_104_2653_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u32_u32_2650_Update/$exit
      -- 
    ca_11138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2650_inst_ack_1, ack => cp_elements(671)); -- 
    rr_11150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(671), ack => EQ_u32_u1_2656_inst_req_0); -- 
    -- CP-element group 672 transition  output  bypass 
    -- predecessors 667 
    -- successors 674 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Update/$entry
      -- 
    cp_elements(672) <= cp_elements(667);
    cr_11155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(672), ack => EQ_u32_u1_2656_inst_req_1); -- 
    -- CP-element group 673 transition  input  bypass 
    -- predecessors 671 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Sample/$exit
      -- 
    ra_11151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2656_inst_ack_0, ack => cp_elements(673)); -- 
    -- CP-element group 674 transition  input  bypass 
    -- predecessors 672 
    -- successors 681 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/EQ_u32_u1_2656_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_105_2667_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_105_2667_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_105_2667_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_105_2667_update_completed_
      -- 
    ca_11156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2656_inst_ack_1, ack => cp_elements(674)); -- 
    -- CP-element group 675 transition  output  bypass 
    -- predecessors 667 
    -- successors 680 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Update/cr
      -- 
    cp_elements(675) <= cp_elements(667);
    cr_11187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(675), ack => NEQ_i32_u1_2664_inst_req_1); -- 
    -- CP-element group 676 transition  output  bypass 
    -- predecessors 667 
    -- successors 677 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2659_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2659_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2659_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_tempx_x0x_xphx_xix_xi_2659_sample_start_
      -- 
    cp_elements(676) <= cp_elements(667);
    rr_11172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(676), ack => type_cast_2660_inst_req_0); -- 
    -- CP-element group 677 transition  input  output  bypass 
    -- predecessors 676 
    -- successors 678 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_sample_completed_
      -- 
    ra_11173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2660_inst_ack_0, ack => cp_elements(677)); -- 
    cr_11177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(677), ack => type_cast_2660_inst_req_1); -- 
    -- CP-element group 678 transition  input  output  bypass 
    -- predecessors 677 
    -- successors 679 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/type_cast_2660_Update/$exit
      -- 
    ca_11178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2660_inst_ack_1, ack => cp_elements(678)); -- 
    rr_11182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => NEQ_i32_u1_2664_inst_req_0); -- 
    -- CP-element group 679 transition  input  bypass 
    -- predecessors 678 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Sample/$exit
      -- 
    ra_11183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2664_inst_ack_0, ack => cp_elements(679)); -- 
    -- CP-element group 680 transition  input  bypass 
    -- predecessors 675 
    -- successors 681 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/NEQ_i32_u1_2664_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_106_2668_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_106_2668_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_106_2668_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/R_iNsTr_106_2668_update_completed_
      -- 
    ca_11188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2664_inst_ack_1, ack => cp_elements(680)); -- 
    -- CP-element group 681 join  transition  output  bypass 
    -- predecessors 674 680 
    -- successors 683 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Sample/rr
      -- 
    cp_element_group_681: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_681"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(674) & cp_elements(680);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(681), clk => clk, reset => reset); --
    end block;
    rr_11204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(681), ack => AND_u1_u1_2669_inst_req_0); -- 
    -- CP-element group 682 transition  output  bypass 
    -- predecessors 667 
    -- successors 684 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Update/cr
      -- 
    cp_elements(682) <= cp_elements(667);
    cr_11209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => AND_u1_u1_2669_inst_req_1); -- 
    -- CP-element group 683 transition  input  bypass 
    -- predecessors 681 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Sample/ra
      -- 
    ra_11205_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2669_inst_ack_0, ack => cp_elements(683)); -- 
    -- CP-element group 684 branch  transition  place  input  bypass 
    -- predecessors 682 
    -- successors 685 686 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2671__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670/AND_u1_u1_2669_Update/ca
      -- 
    ca_11210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2669_inst_ack_1, ack => cp_elements(684)); -- 
    -- CP-element group 685 transition  place  dead  bypass 
    -- predecessors 684 
    -- successors 38 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2677__entry__
      -- 	branch_block_stmt_1659/if_stmt_2671__exit__
      -- 	branch_block_stmt_1659/if_stmt_2671_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2671_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2671_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2677_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2677_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2677_dead_link/dead_transition
      -- 
    cp_elements(685) <= false;
    -- CP-element group 686 transition  output  bypass 
    -- predecessors 684 
    -- successors 687 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2671_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2671_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2671_eval_test/branch_req
      -- 
    cp_elements(686) <= cp_elements(684);
    branch_req_11218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => if_stmt_2671_branch_req_0); -- 
    -- CP-element group 687 branch  place  bypass 
    -- predecessors 686 
    -- successors 688 690 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcond11x_xix_xi_2672_place
      -- 
    cp_elements(687) <= cp_elements(686);
    -- CP-element group 688 transition  bypass 
    -- predecessors 687 
    -- successors 689 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2671_if_link/$entry
      -- 
    cp_elements(688) <= cp_elements(687);
    -- CP-element group 689 transition  place  input  bypass 
    -- predecessors 688 
    -- successors 38 
    -- members (9) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader
      -- 	branch_block_stmt_1659/if_stmt_2671_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2671_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_udiv32x_xexitx_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2677_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_2677_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2677_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2677_PhiAck/dummy
      -- 
    if_choice_transition_11223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2671_branch_ack_1, ack => cp_elements(689)); -- 
    -- CP-element group 690 transition  bypass 
    -- predecessors 687 
    -- successors 691 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2671_else_link/$entry
      -- 
    cp_elements(690) <= cp_elements(687);
    -- CP-element group 691 transition  place  input  bypass 
    -- predecessors 690 
    -- successors 1818 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_2671_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2671_else_link/else_choice_transition
      -- 
    else_choice_transition_11227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2671_branch_ack_0, ack => cp_elements(691)); -- 
    -- CP-element group 692 fork  transition  bypass 
    -- predecessors 39 
    -- successors 693 694 697 701 704 711 714 715 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/$entry
      -- 
    cp_elements(692) <= cp_elements(39);
    -- CP-element group 693 transition  output  bypass 
    -- predecessors 692 
    -- successors 696 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Update/cr
      -- 
    cp_elements(693) <= cp_elements(692);
    cr_11249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => SHL_u32_u32_2698_inst_req_1); -- 
    -- CP-element group 694 transition  output  bypass 
    -- predecessors 692 
    -- successors 695 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_tempx_x012x_xix_xi_2695_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_tempx_x012x_xix_xi_2695_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_tempx_x012x_xix_xi_2695_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_tempx_x012x_xix_xi_2695_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Sample/rr
      -- 
    cp_elements(694) <= cp_elements(692);
    rr_11244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => SHL_u32_u32_2698_inst_req_0); -- 
    -- CP-element group 695 transition  input  bypass 
    -- predecessors 694 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Sample/ra
      -- 
    ra_11245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2698_inst_ack_0, ack => cp_elements(695)); -- 
    -- CP-element group 696 fork  transition  input  bypass 
    -- predecessors 693 
    -- successors 698 705 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/SHL_u32_u32_2698_Update/ca
      -- 
    ca_11250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2698_inst_ack_1, ack => cp_elements(696)); -- 
    -- CP-element group 697 transition  output  bypass 
    -- predecessors 692 
    -- successors 700 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Update/cr
      -- 
    cp_elements(697) <= cp_elements(692);
    cr_11267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => AND_u32_u32_2704_inst_req_1); -- 
    -- CP-element group 698 transition  output  bypass 
    -- predecessors 696 
    -- successors 699 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2701_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2701_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2701_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2701_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Sample/rr
      -- 
    cp_elements(698) <= cp_elements(696);
    rr_11262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(698), ack => AND_u32_u32_2704_inst_req_0); -- 
    -- CP-element group 699 transition  input  bypass 
    -- predecessors 698 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Sample/ra
      -- 
    ra_11263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2704_inst_ack_0, ack => cp_elements(699)); -- 
    -- CP-element group 700 transition  input  output  bypass 
    -- predecessors 697 
    -- successors 702 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u32_u32_2704_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_158_2707_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_158_2707_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_158_2707_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_158_2707_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Sample/rr
      -- 
    ca_11268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2704_inst_ack_1, ack => cp_elements(700)); -- 
    rr_11280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(700), ack => EQ_u32_u1_2710_inst_req_0); -- 
    -- CP-element group 701 transition  output  bypass 
    -- predecessors 692 
    -- successors 703 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Update/cr
      -- 
    cp_elements(701) <= cp_elements(692);
    cr_11285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => EQ_u32_u1_2710_inst_req_1); -- 
    -- CP-element group 702 transition  input  bypass 
    -- predecessors 700 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Sample/ra
      -- 
    ra_11281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2710_inst_ack_0, ack => cp_elements(702)); -- 
    -- CP-element group 703 transition  input  bypass 
    -- predecessors 701 
    -- successors 710 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/EQ_u32_u1_2710_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_159_2721_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_159_2721_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_159_2721_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_159_2721_update_completed_
      -- 
    ca_11286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2710_inst_ack_1, ack => cp_elements(703)); -- 
    -- CP-element group 704 transition  output  bypass 
    -- predecessors 692 
    -- successors 709 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Update/cr
      -- 
    cp_elements(704) <= cp_elements(692);
    cr_11317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(704), ack => NEQ_i32_u1_2718_inst_req_1); -- 
    -- CP-element group 705 transition  output  bypass 
    -- predecessors 696 
    -- successors 706 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2713_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2713_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2713_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_157_2713_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Sample/rr
      -- 
    cp_elements(705) <= cp_elements(696);
    rr_11302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => type_cast_2714_inst_req_0); -- 
    -- CP-element group 706 transition  input  output  bypass 
    -- predecessors 705 
    -- successors 707 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Update/cr
      -- 
    ra_11303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_0, ack => cp_elements(706)); -- 
    cr_11307_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(706), ack => type_cast_2714_inst_req_1); -- 
    -- CP-element group 707 transition  input  output  bypass 
    -- predecessors 706 
    -- successors 708 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/type_cast_2714_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Sample/rr
      -- 
    ca_11308_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_1, ack => cp_elements(707)); -- 
    rr_11312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => NEQ_i32_u1_2718_inst_req_0); -- 
    -- CP-element group 708 transition  input  bypass 
    -- predecessors 707 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Sample/ra
      -- 
    ra_11313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2718_inst_ack_0, ack => cp_elements(708)); -- 
    -- CP-element group 709 transition  input  bypass 
    -- predecessors 704 
    -- successors 710 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/NEQ_i32_u1_2718_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_160_2722_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_160_2722_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_160_2722_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_160_2722_update_completed_
      -- 
    ca_11318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_2718_inst_ack_1, ack => cp_elements(709)); -- 
    -- CP-element group 710 join  transition  output  bypass 
    -- predecessors 703 709 
    -- successors 712 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Sample/rr
      -- 
    cp_element_group_710: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_710"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(703) & cp_elements(709);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(710), clk => clk, reset => reset); --
    end block;
    rr_11334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => AND_u1_u1_2723_inst_req_0); -- 
    -- CP-element group 711 transition  output  bypass 
    -- predecessors 692 
    -- successors 713 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Update/cr
      -- 
    cp_elements(711) <= cp_elements(692);
    cr_11339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => AND_u1_u1_2723_inst_req_1); -- 
    -- CP-element group 712 transition  input  bypass 
    -- predecessors 710 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Sample/ra
      -- 
    ra_11335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2723_inst_ack_0, ack => cp_elements(712)); -- 
    -- CP-element group 713 transition  input  bypass 
    -- predecessors 711 
    -- successors 718 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/AND_u1_u1_2723_Update/ca
      -- 
    ca_11340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2723_inst_ack_1, ack => cp_elements(713)); -- 
    -- CP-element group 714 transition  output  bypass 
    -- predecessors 692 
    -- successors 717 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Update/cr
      -- 
    cp_elements(714) <= cp_elements(692);
    cr_11357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(714), ack => ADD_u32_u32_2729_inst_req_1); -- 
    -- CP-element group 715 transition  output  bypass 
    -- predecessors 692 
    -- successors 716 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_156_2726_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_156_2726_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_156_2726_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/R_iNsTr_156_2726_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Sample/rr
      -- 
    cp_elements(715) <= cp_elements(692);
    rr_11352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(715), ack => ADD_u32_u32_2729_inst_req_0); -- 
    -- CP-element group 716 transition  input  bypass 
    -- predecessors 715 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Sample/ra
      -- 
    ra_11353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2729_inst_ack_0, ack => cp_elements(716)); -- 
    -- CP-element group 717 transition  input  bypass 
    -- predecessors 714 
    -- successors 718 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/ADD_u32_u32_2729_Update/ca
      -- 
    ca_11358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2729_inst_ack_1, ack => cp_elements(717)); -- 
    -- CP-element group 718 join  transition  bypass 
    -- predecessors 713 717 
    -- successors 40 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2699_to_assign_stmt_2730/$exit
      -- 
    cp_element_group_718: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_718"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(713) & cp_elements(717);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(718), clk => clk, reset => reset); --
    end block;
    -- CP-element group 719 transition  place  dead  bypass 
    -- predecessors 40 
    -- successors 41 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2737__entry__
      -- 	branch_block_stmt_1659/if_stmt_2731__exit__
      -- 	branch_block_stmt_1659/if_stmt_2731_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2731_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2731_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2737_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2737_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2737_dead_link/dead_transition
      -- 
    cp_elements(719) <= false;
    -- CP-element group 720 transition  output  bypass 
    -- predecessors 40 
    -- successors 721 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2731_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2731_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2731_eval_test/branch_req
      -- 
    cp_elements(720) <= cp_elements(40);
    branch_req_11366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => if_stmt_2731_branch_req_0); -- 
    -- CP-element group 721 branch  place  bypass 
    -- predecessors 720 
    -- successors 722 724 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcondx_xix_xi_2732_place
      -- 
    cp_elements(721) <= cp_elements(720);
    -- CP-element group 722 transition  bypass 
    -- predecessors 721 
    -- successors 723 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2731_if_link/$entry
      -- 
    cp_elements(722) <= cp_elements(721);
    -- CP-element group 723 transition  place  input  bypass 
    -- predecessors 722 
    -- successors 1756 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_2731_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2731_if_link/if_choice_transition
      -- 
    if_choice_transition_11371_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2731_branch_ack_1, ack => cp_elements(723)); -- 
    -- CP-element group 724 transition  bypass 
    -- predecessors 721 
    -- successors 725 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2731_else_link/$entry
      -- 
    cp_elements(724) <= cp_elements(721);
    -- CP-element group 725 transition  place  input  bypass 
    -- predecessors 724 
    -- successors 1799 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_2731_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2731_else_link/else_choice_transition
      -- 
    else_choice_transition_11375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2731_branch_ack_0, ack => cp_elements(725)); -- 
    -- CP-element group 726 fork  transition  bypass 
    -- predecessors 41 
    -- successors 727 728 731 735 736 740 741 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/$entry
      -- 
    cp_elements(726) <= cp_elements(41);
    -- CP-element group 727 transition  output  bypass 
    -- predecessors 726 
    -- successors 730 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Update/cr
      -- 
    cp_elements(727) <= cp_elements(726);
    cr_11397_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => OR_u32_u32_2751_inst_req_1); -- 
    -- CP-element group 728 transition  output  bypass 
    -- predecessors 726 
    -- successors 729 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_78_2748_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_78_2748_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_78_2748_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_78_2748_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Sample/rr
      -- 
    cp_elements(728) <= cp_elements(726);
    rr_11392_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => OR_u32_u32_2751_inst_req_0); -- 
    -- CP-element group 729 transition  input  bypass 
    -- predecessors 728 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Sample/ra
      -- 
    ra_11393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2751_inst_ack_0, ack => cp_elements(729)); -- 
    -- CP-element group 730 transition  input  output  bypass 
    -- predecessors 727 
    -- successors 732 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/OR_u32_u32_2751_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xnotx_xi_2754_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xnotx_xi_2754_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xnotx_xi_2754_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xnotx_xi_2754_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Sample/rr
      -- 
    ca_11398_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2751_inst_ack_1, ack => cp_elements(730)); -- 
    rr_11410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(730), ack => XOR_u32_u32_2757_inst_req_0); -- 
    -- CP-element group 731 transition  output  bypass 
    -- predecessors 726 
    -- successors 733 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Update/cr
      -- 
    cp_elements(731) <= cp_elements(726);
    cr_11415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(731), ack => XOR_u32_u32_2757_inst_req_1); -- 
    -- CP-element group 732 transition  input  bypass 
    -- predecessors 730 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Sample/ra
      -- 
    ra_11411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2757_inst_ack_0, ack => cp_elements(732)); -- 
    -- CP-element group 733 transition  input  bypass 
    -- predecessors 731 
    -- successors 734 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/XOR_u32_u32_2757_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp21x_xix_xi_2761_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp21x_xix_xi_2761_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp21x_xix_xi_2761_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp21x_xix_xi_2761_update_completed_
      -- 
    ca_11416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_2757_inst_ack_1, ack => cp_elements(733)); -- 
    -- CP-element group 734 join  transition  output  bypass 
    -- predecessors 733 736 
    -- successors 737 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Sample/rr
      -- 
    cp_element_group_734: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_734"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(733) & cp_elements(736);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(734), clk => clk, reset => reset); --
    end block;
    rr_11432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => ADD_u32_u32_2762_inst_req_0); -- 
    -- CP-element group 735 transition  output  bypass 
    -- predecessors 726 
    -- successors 738 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Update/cr
      -- 
    cp_elements(735) <= cp_elements(726);
    cr_11437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => ADD_u32_u32_2762_inst_req_1); -- 
    -- CP-element group 736 transition  bypass 
    -- predecessors 726 
    -- successors 734 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_77_2760_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_77_2760_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_77_2760_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_iNsTr_77_2760_update_completed_
      -- 
    cp_elements(736) <= cp_elements(726);
    -- CP-element group 737 transition  input  bypass 
    -- predecessors 734 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Sample/ra
      -- 
    ra_11433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2762_inst_ack_0, ack => cp_elements(737)); -- 
    -- CP-element group 738 transition  input  bypass 
    -- predecessors 735 
    -- successors 739 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/ADD_u32_u32_2762_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp25x_xix_xi_2765_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp25x_xix_xi_2765_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp25x_xix_xi_2765_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_tmp25x_xix_xi_2765_update_completed_
      -- 
    ca_11438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2762_inst_ack_1, ack => cp_elements(738)); -- 
    -- CP-element group 739 join  transition  output  bypass 
    -- predecessors 738 741 
    -- successors 742 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Sample/rr
      -- 
    cp_element_group_739: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_739"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(738) & cp_elements(741);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(739), clk => clk, reset => reset); --
    end block;
    rr_11454_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => SUB_u32_u32_2767_inst_req_0); -- 
    -- CP-element group 740 transition  output  bypass 
    -- predecessors 726 
    -- successors 743 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Update/cr
      -- 
    cp_elements(740) <= cp_elements(726);
    cr_11459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => SUB_u32_u32_2767_inst_req_1); -- 
    -- CP-element group 741 transition  bypass 
    -- predecessors 726 
    -- successors 739 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xlcssa5_2766_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xlcssa5_2766_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xlcssa5_2766_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/R_xx_xlcssa5_2766_update_completed_
      -- 
    cp_elements(741) <= cp_elements(726);
    -- CP-element group 742 transition  input  bypass 
    -- predecessors 739 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Sample/ra
      -- 
    ra_11455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2767_inst_ack_0, ack => cp_elements(742)); -- 
    -- CP-element group 743 transition  place  input  bypass 
    -- predecessors 740 
    -- successors 1844 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768__exit__
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2752_to_assign_stmt_2768/SUB_u32_u32_2767_Update/ca
      -- 
    ca_11460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_2767_inst_ack_1, ack => cp_elements(743)); -- 
    -- CP-element group 744 fork  transition  bypass 
    -- predecessors 42 
    -- successors 745 746 749 750 753 757 758 762 765 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/$entry
      -- 
    cp_elements(744) <= cp_elements(42);
    -- CP-element group 745 transition  output  bypass 
    -- predecessors 744 
    -- successors 748 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Update/cr
      -- 
    cp_elements(745) <= cp_elements(744);
    cr_11480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => AND_u32_u32_2788_inst_req_1); -- 
    -- CP-element group 746 transition  output  bypass 
    -- predecessors 744 
    -- successors 747 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_tempx_x0x_xlcssax_xix_xi_2785_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_tempx_x0x_xlcssax_xix_xi_2785_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_tempx_x0x_xlcssax_xix_xi_2785_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_tempx_x0x_xlcssax_xix_xi_2785_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Sample/rr
      -- 
    cp_elements(746) <= cp_elements(744);
    rr_11475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(746), ack => AND_u32_u32_2788_inst_req_0); -- 
    -- CP-element group 747 transition  input  bypass 
    -- predecessors 746 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Sample/ra
      -- 
    ra_11476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2788_inst_ack_0, ack => cp_elements(747)); -- 
    -- CP-element group 748 transition  input  bypass 
    -- predecessors 745 
    -- successors 756 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/AND_u32_u32_2788_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_129_2803_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_129_2803_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_129_2803_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_129_2803_update_completed_
      -- 
    ca_11481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2788_inst_ack_1, ack => cp_elements(748)); -- 
    -- CP-element group 749 transition  output  bypass 
    -- predecessors 744 
    -- successors 752 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Update/cr
      -- 
    cp_elements(749) <= cp_elements(744);
    cr_11498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => SHL_u32_u32_2794_inst_req_1); -- 
    -- CP-element group 750 transition  output  bypass 
    -- predecessors 744 
    -- successors 751 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_expx_x0x_xlcssax_xix_xi_2791_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_expx_x0x_xlcssax_xix_xi_2791_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_expx_x0x_xlcssax_xix_xi_2791_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_expx_x0x_xlcssax_xix_xi_2791_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Sample/rr
      -- 
    cp_elements(750) <= cp_elements(744);
    rr_11493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(750), ack => SHL_u32_u32_2794_inst_req_0); -- 
    -- CP-element group 751 transition  input  bypass 
    -- predecessors 750 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Sample/ra
      -- 
    ra_11494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2794_inst_ack_0, ack => cp_elements(751)); -- 
    -- CP-element group 752 transition  input  output  bypass 
    -- predecessors 749 
    -- successors 754 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/SHL_u32_u32_2794_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_130_2797_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_130_2797_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_130_2797_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_130_2797_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Sample/rr
      -- 
    ca_11499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2794_inst_ack_1, ack => cp_elements(752)); -- 
    rr_11511_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(752), ack => ADD_u32_u32_2800_inst_req_0); -- 
    -- CP-element group 753 transition  output  bypass 
    -- predecessors 744 
    -- successors 755 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Update/cr
      -- 
    cp_elements(753) <= cp_elements(744);
    cr_11516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ADD_u32_u32_2800_inst_req_1); -- 
    -- CP-element group 754 transition  input  bypass 
    -- predecessors 752 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Sample/ra
      -- 
    ra_11512_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2800_inst_ack_0, ack => cp_elements(754)); -- 
    -- CP-element group 755 transition  input  bypass 
    -- predecessors 753 
    -- successors 761 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/ADD_u32_u32_2800_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_131_2809_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_131_2809_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_131_2809_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_131_2809_update_completed_
      -- 
    ca_11517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2800_inst_ack_1, ack => cp_elements(755)); -- 
    -- CP-element group 756 join  transition  output  bypass 
    -- predecessors 748 758 
    -- successors 759 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Sample/rr
      -- 
    cp_element_group_756: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_756"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(748) & cp_elements(758);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(756), clk => clk, reset => reset); --
    end block;
    rr_11533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => OR_u32_u32_2805_inst_req_0); -- 
    -- CP-element group 757 transition  output  bypass 
    -- predecessors 744 
    -- successors 760 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Update/cr
      -- 
    cp_elements(757) <= cp_elements(744);
    cr_11538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => OR_u32_u32_2805_inst_req_1); -- 
    -- CP-element group 758 transition  bypass 
    -- predecessors 744 
    -- successors 756 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_87_2804_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_87_2804_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_87_2804_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_87_2804_update_completed_
      -- 
    cp_elements(758) <= cp_elements(744);
    -- CP-element group 759 transition  input  bypass 
    -- predecessors 756 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Sample/ra
      -- 
    ra_11534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2805_inst_ack_0, ack => cp_elements(759)); -- 
    -- CP-element group 760 transition  input  bypass 
    -- predecessors 757 
    -- successors 761 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2805_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_132_2808_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_132_2808_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_132_2808_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_132_2808_update_completed_
      -- 
    ca_11539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2805_inst_ack_1, ack => cp_elements(760)); -- 
    -- CP-element group 761 join  transition  output  bypass 
    -- predecessors 755 760 
    -- successors 763 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Sample/rr
      -- 
    cp_element_group_761: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_761"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(755) & cp_elements(760);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(761), clk => clk, reset => reset); --
    end block;
    rr_11555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => OR_u32_u32_2810_inst_req_0); -- 
    -- CP-element group 762 transition  output  bypass 
    -- predecessors 744 
    -- successors 764 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Update/cr
      -- 
    cp_elements(762) <= cp_elements(744);
    cr_11560_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(762), ack => OR_u32_u32_2810_inst_req_1); -- 
    -- CP-element group 763 transition  input  bypass 
    -- predecessors 761 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Sample/ra
      -- 
    ra_11556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2810_inst_ack_0, ack => cp_elements(763)); -- 
    -- CP-element group 764 transition  input  output  bypass 
    -- predecessors 762 
    -- successors 766 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/OR_u32_u32_2810_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_133_2813_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_133_2813_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_133_2813_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/R_iNsTr_133_2813_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Sample/rr
      -- 
    ca_11561_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2810_inst_ack_1, ack => cp_elements(764)); -- 
    rr_11573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(764), ack => type_cast_2814_inst_req_0); -- 
    -- CP-element group 765 transition  output  bypass 
    -- predecessors 744 
    -- successors 767 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Update/cr
      -- 
    cp_elements(765) <= cp_elements(744);
    cr_11578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => type_cast_2814_inst_req_1); -- 
    -- CP-element group 766 transition  input  bypass 
    -- predecessors 764 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Sample/ra
      -- 
    ra_11574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2814_inst_ack_0, ack => cp_elements(766)); -- 
    -- CP-element group 767 fork  transition  place  input  bypass 
    -- predecessors 765 
    -- successors 1878 1880 
    -- members (11) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2789_to_assign_stmt_2815/type_cast_2814_Update/ca
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/$entry
      -- 
    ca_11579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2814_inst_ack_1, ack => cp_elements(767)); -- 
    -- CP-element group 768 fork  transition  bypass 
    -- predecessors 1885 
    -- successors 769 770 774 775 778 781 785 786 789 792 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/$entry
      -- 
    cp_elements(768) <= cp_elements(1885);
    -- CP-element group 769 transition  output  bypass 
    -- predecessors 768 
    -- successors 772 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Update/cr
      -- 
    cp_elements(769) <= cp_elements(768);
    cr_11599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(769), ack => MUL_f32_f32_2830_inst_req_1); -- 
    -- CP-element group 770 transition  output  bypass 
    -- predecessors 768 
    -- successors 771 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_39_2827_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_39_2827_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_39_2827_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_39_2827_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Sample/rr
      -- 
    cp_elements(770) <= cp_elements(768);
    rr_11594_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => MUL_f32_f32_2830_inst_req_0); -- 
    -- CP-element group 771 transition  input  bypass 
    -- predecessors 770 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Sample/ra
      -- 
    ra_11595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2830_inst_ack_0, ack => cp_elements(771)); -- 
    -- CP-element group 772 transition  input  bypass 
    -- predecessors 769 
    -- successors 773 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2830_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_68_2833_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_68_2833_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_68_2833_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_68_2833_update_completed_
      -- 
    ca_11600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2830_inst_ack_1, ack => cp_elements(772)); -- 
    -- CP-element group 773 join  transition  output  bypass 
    -- predecessors 772 775 
    -- successors 776 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Sample/rr
      -- 
    cp_element_group_773: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_773"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(772) & cp_elements(775);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(773), clk => clk, reset => reset); --
    end block;
    rr_11616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(773), ack => ADD_f32_f32_2835_inst_req_0); -- 
    -- CP-element group 774 transition  output  bypass 
    -- predecessors 768 
    -- successors 777 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Update/cr
      -- 
    cp_elements(774) <= cp_elements(768);
    cr_11621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => ADD_f32_f32_2835_inst_req_1); -- 
    -- CP-element group 775 transition  bypass 
    -- predecessors 768 
    -- successors 773 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_flux_rotor_lpf_prevx_x0_2834_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_flux_rotor_lpf_prevx_x0_2834_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_flux_rotor_lpf_prevx_x0_2834_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_flux_rotor_lpf_prevx_x0_2834_update_completed_
      -- 
    cp_elements(775) <= cp_elements(768);
    -- CP-element group 776 transition  input  bypass 
    -- predecessors 773 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Sample/ra
      -- 
    ra_11617_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2835_inst_ack_0, ack => cp_elements(776)); -- 
    -- CP-element group 777 transition  input  output  bypass 
    -- predecessors 774 
    -- successors 779 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2835_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_69_2840_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_69_2840_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_69_2840_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_69_2840_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Sample/rr
      -- 
    ca_11622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2835_inst_ack_1, ack => cp_elements(777)); -- 
    rr_11634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(777), ack => SUB_f32_f32_2841_inst_req_0); -- 
    -- CP-element group 778 transition  output  bypass 
    -- predecessors 768 
    -- successors 780 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Update/cr
      -- 
    cp_elements(778) <= cp_elements(768);
    cr_11639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(778), ack => SUB_f32_f32_2841_inst_req_1); -- 
    -- CP-element group 779 transition  input  bypass 
    -- predecessors 777 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Sample/ra
      -- 
    ra_11635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2841_inst_ack_0, ack => cp_elements(779)); -- 
    -- CP-element group 780 transition  input  output  bypass 
    -- predecessors 778 
    -- successors 782 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SUB_f32_f32_2841_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_70_2844_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_70_2844_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_70_2844_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_70_2844_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Sample/rr
      -- 
    ca_11640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2841_inst_ack_1, ack => cp_elements(780)); -- 
    rr_11652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(780), ack => MUL_f32_f32_2847_inst_req_0); -- 
    -- CP-element group 781 transition  output  bypass 
    -- predecessors 768 
    -- successors 783 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Update/cr
      -- 
    cp_elements(781) <= cp_elements(768);
    cr_11657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(781), ack => MUL_f32_f32_2847_inst_req_1); -- 
    -- CP-element group 782 transition  input  bypass 
    -- predecessors 780 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Sample/ra
      -- 
    ra_11653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2847_inst_ack_0, ack => cp_elements(782)); -- 
    -- CP-element group 783 transition  input  bypass 
    -- predecessors 781 
    -- successors 784 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2847_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_71_2850_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_71_2850_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_71_2850_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_71_2850_update_completed_
      -- 
    ca_11658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2847_inst_ack_1, ack => cp_elements(783)); -- 
    -- CP-element group 784 join  transition  output  bypass 
    -- predecessors 783 786 
    -- successors 787 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Sample/rr
      -- 
    cp_element_group_784: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_784"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(783) & cp_elements(786);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(784), clk => clk, reset => reset); --
    end block;
    rr_11674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => ADD_f32_f32_2852_inst_req_0); -- 
    -- CP-element group 785 transition  output  bypass 
    -- predecessors 768 
    -- successors 788 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Update/cr
      -- 
    cp_elements(785) <= cp_elements(768);
    cr_11679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => ADD_f32_f32_2852_inst_req_1); -- 
    -- CP-element group 786 transition  bypass 
    -- predecessors 768 
    -- successors 784 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_int_flux_err_temp_2x_x0_2851_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_int_flux_err_temp_2x_x0_2851_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_int_flux_err_temp_2x_x0_2851_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_int_flux_err_temp_2x_x0_2851_update_completed_
      -- 
    cp_elements(786) <= cp_elements(768);
    -- CP-element group 787 transition  input  bypass 
    -- predecessors 784 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Sample/ra
      -- 
    ra_11675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2852_inst_ack_0, ack => cp_elements(787)); -- 
    -- CP-element group 788 transition  input  output  bypass 
    -- predecessors 785 
    -- successors 790 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/ADD_f32_f32_2852_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_72_2855_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_72_2855_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_72_2855_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_72_2855_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Sample/rr
      -- 
    ca_11680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2852_inst_ack_1, ack => cp_elements(788)); -- 
    rr_11692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => MUL_f32_f32_2858_inst_req_0); -- 
    -- CP-element group 789 transition  output  bypass 
    -- predecessors 768 
    -- successors 791 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Update/cr
      -- 
    cp_elements(789) <= cp_elements(768);
    cr_11697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(789), ack => MUL_f32_f32_2858_inst_req_1); -- 
    -- CP-element group 790 transition  input  bypass 
    -- predecessors 788 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Sample/ra
      -- 
    ra_11693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2858_inst_ack_0, ack => cp_elements(790)); -- 
    -- CP-element group 791 transition  input  output  bypass 
    -- predecessors 789 
    -- successors 793 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/MUL_f32_f32_2858_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_73_2861_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_73_2861_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_73_2861_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/R_iNsTr_73_2861_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Sample/rr
      -- 
    ca_11698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2858_inst_ack_1, ack => cp_elements(791)); -- 
    rr_11710_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => SLT_f32_u1_2864_inst_req_0); -- 
    -- CP-element group 792 transition  output  bypass 
    -- predecessors 768 
    -- successors 794 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Update/cr
      -- 
    cp_elements(792) <= cp_elements(768);
    cr_11715_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(792), ack => SLT_f32_u1_2864_inst_req_1); -- 
    -- CP-element group 793 transition  input  bypass 
    -- predecessors 791 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Sample/ra
      -- 
    ra_11711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2864_inst_ack_0, ack => cp_elements(793)); -- 
    -- CP-element group 794 branch  transition  place  input  bypass 
    -- predecessors 792 
    -- successors 795 796 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2866__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865/SLT_f32_u1_2864_Update/ca
      -- 
    ca_11716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2864_inst_ack_1, ack => cp_elements(794)); -- 
    -- CP-element group 795 transition  place  dead  bypass 
    -- predecessors 794 
    -- successors 43 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2872__entry__
      -- 	branch_block_stmt_1659/if_stmt_2866__exit__
      -- 	branch_block_stmt_1659/if_stmt_2866_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2866_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2866_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2872_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2872_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2872_dead_link/$entry
      -- 
    cp_elements(795) <= false;
    -- CP-element group 796 transition  output  bypass 
    -- predecessors 794 
    -- successors 797 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2866_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2866_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2866_eval_test/branch_req
      -- 
    cp_elements(796) <= cp_elements(794);
    branch_req_11724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => if_stmt_2866_branch_req_0); -- 
    -- CP-element group 797 branch  place  bypass 
    -- predecessors 796 
    -- successors 798 800 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_74_2867_place
      -- 
    cp_elements(797) <= cp_elements(796);
    -- CP-element group 798 transition  bypass 
    -- predecessors 797 
    -- successors 799 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2866_if_link/$entry
      -- 
    cp_elements(798) <= cp_elements(797);
    -- CP-element group 799 fork  transition  place  input  bypass 
    -- predecessors 798 
    -- successors 1894 1895 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2866_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2866_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$entry
      -- 
    if_choice_transition_11729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2866_branch_ack_1, ack => cp_elements(799)); -- 
    -- CP-element group 800 transition  bypass 
    -- predecessors 797 
    -- successors 801 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2866_else_link/$entry
      -- 
    cp_elements(800) <= cp_elements(797);
    -- CP-element group 801 transition  place  input  bypass 
    -- predecessors 800 
    -- successors 43 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2866_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2866_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_42
      -- 	branch_block_stmt_1659/merge_stmt_2872_PhiAck/dummy
      -- 	branch_block_stmt_1659/merge_stmt_2872_PhiAck/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_42_PhiReq/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_42_PhiReq/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2872_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2872_PhiReqMerge
      -- 
    else_choice_transition_11733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2866_branch_ack_0, ack => cp_elements(801)); -- 
    -- CP-element group 802 fork  transition  bypass 
    -- predecessors 43 
    -- successors 803 804 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2878/$entry
      -- 
    cp_elements(802) <= cp_elements(43);
    -- CP-element group 803 transition  output  bypass 
    -- predecessors 802 
    -- successors 806 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Update/cr
      -- 
    cp_elements(803) <= cp_elements(802);
    cr_11755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => SGT_f32_u1_2877_inst_req_1); -- 
    -- CP-element group 804 transition  output  bypass 
    -- predecessors 802 
    -- successors 805 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2878/R_iNsTr_73_2874_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2878/R_iNsTr_73_2874_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2878/R_iNsTr_73_2874_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2878/R_iNsTr_73_2874_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Sample/rr
      -- 
    cp_elements(804) <= cp_elements(802);
    rr_11750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => SGT_f32_u1_2877_inst_req_0); -- 
    -- CP-element group 805 transition  input  bypass 
    -- predecessors 804 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Sample/ra
      -- 
    ra_11751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2877_inst_ack_0, ack => cp_elements(805)); -- 
    -- CP-element group 806 branch  transition  place  input  bypass 
    -- predecessors 803 
    -- successors 807 808 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2879__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2878__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2878/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2878/SGT_f32_u1_2877_Update/ca
      -- 
    ca_11756_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2877_inst_ack_1, ack => cp_elements(806)); -- 
    -- CP-element group 807 transition  place  dead  bypass 
    -- predecessors 806 
    -- successors 44 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2885__entry__
      -- 	branch_block_stmt_1659/if_stmt_2879__exit__
      -- 	branch_block_stmt_1659/if_stmt_2879_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2879_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2879_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2885_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2885_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2885_dead_link/dead_transition
      -- 
    cp_elements(807) <= false;
    -- CP-element group 808 transition  output  bypass 
    -- predecessors 806 
    -- successors 809 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2879_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2879_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2879_eval_test/branch_req
      -- 
    cp_elements(808) <= cp_elements(806);
    branch_req_11764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => if_stmt_2879_branch_req_0); -- 
    -- CP-element group 809 branch  place  bypass 
    -- predecessors 808 
    -- successors 810 812 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_100_2880_place
      -- 
    cp_elements(809) <= cp_elements(808);
    -- CP-element group 810 transition  bypass 
    -- predecessors 809 
    -- successors 811 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2879_if_link/$entry
      -- 
    cp_elements(810) <= cp_elements(809);
    -- CP-element group 811 fork  transition  place  input  bypass 
    -- predecessors 810 
    -- successors 1886 1887 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2879_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2879_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_42_bb_44
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$entry
      -- 
    if_choice_transition_11769_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2879_branch_ack_1, ack => cp_elements(811)); -- 
    -- CP-element group 812 transition  bypass 
    -- predecessors 809 
    -- successors 813 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2879_else_link/$entry
      -- 
    cp_elements(812) <= cp_elements(809);
    -- CP-element group 813 transition  place  input  bypass 
    -- predecessors 812 
    -- successors 44 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2879_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2879_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_42_bb_43
      -- 	branch_block_stmt_1659/bb_42_bb_43_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_43_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2885_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2885_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2885_PhiAck/dummy
      -- 	branch_block_stmt_1659/merge_stmt_2885_PhiReqMerge
      -- 
    else_choice_transition_11773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2879_branch_ack_0, ack => cp_elements(813)); -- 
    -- CP-element group 814 fork  transition  bypass 
    -- predecessors 1899 
    -- successors 815 816 820 821 824 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/$entry
      -- 
    cp_elements(814) <= cp_elements(1899);
    -- CP-element group 815 transition  output  bypass 
    -- predecessors 814 
    -- successors 818 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Update/cr
      -- 
    cp_elements(815) <= cp_elements(814);
    cr_11795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => MUL_f32_f32_2903_inst_req_1); -- 
    -- CP-element group 816 transition  output  bypass 
    -- predecessors 814 
    -- successors 817 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_70_2900_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_70_2900_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_70_2900_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_70_2900_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Sample/rr
      -- 
    cp_elements(816) <= cp_elements(814);
    rr_11790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(816), ack => MUL_f32_f32_2903_inst_req_0); -- 
    -- CP-element group 817 transition  input  bypass 
    -- predecessors 816 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Sample/ra
      -- 
    ra_11791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2903_inst_ack_0, ack => cp_elements(817)); -- 
    -- CP-element group 818 transition  input  bypass 
    -- predecessors 815 
    -- successors 819 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/MUL_f32_f32_2903_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_96_2907_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_96_2907_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_96_2907_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_96_2907_update_completed_
      -- 
    ca_11796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_2903_inst_ack_1, ack => cp_elements(818)); -- 
    -- CP-element group 819 join  transition  output  bypass 
    -- predecessors 818 821 
    -- successors 822 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Sample/rr
      -- 
    cp_element_group_819: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_819"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(818) & cp_elements(821);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(819), clk => clk, reset => reset); --
    end block;
    rr_11812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => ADD_f32_f32_2908_inst_req_0); -- 
    -- CP-element group 820 transition  output  bypass 
    -- predecessors 814 
    -- successors 823 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Update/cr
      -- 
    cp_elements(820) <= cp_elements(814);
    cr_11817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(820), ack => ADD_f32_f32_2908_inst_req_1); -- 
    -- CP-element group 821 transition  bypass 
    -- predecessors 814 
    -- successors 819 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_int_flux_errx_x0_2906_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_int_flux_errx_x0_2906_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_int_flux_errx_x0_2906_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_int_flux_errx_x0_2906_update_completed_
      -- 
    cp_elements(821) <= cp_elements(814);
    -- CP-element group 822 transition  input  bypass 
    -- predecessors 819 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Sample/ra
      -- 
    ra_11813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2908_inst_ack_0, ack => cp_elements(822)); -- 
    -- CP-element group 823 transition  input  output  bypass 
    -- predecessors 820 
    -- successors 825 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/ADD_f32_f32_2908_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_97_2911_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_97_2911_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_97_2911_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/R_iNsTr_97_2911_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Sample/rr
      -- 
    ca_11818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2908_inst_ack_1, ack => cp_elements(823)); -- 
    rr_11830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => SLT_f32_u1_2914_inst_req_0); -- 
    -- CP-element group 824 transition  output  bypass 
    -- predecessors 814 
    -- successors 826 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Update/cr
      -- 
    cp_elements(824) <= cp_elements(814);
    cr_11835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(824), ack => SLT_f32_u1_2914_inst_req_1); -- 
    -- CP-element group 825 transition  input  bypass 
    -- predecessors 823 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Sample/ra
      -- 
    ra_11831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2914_inst_ack_0, ack => cp_elements(825)); -- 
    -- CP-element group 826 branch  transition  place  input  bypass 
    -- predecessors 824 
    -- successors 827 828 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2916__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915/SLT_f32_u1_2914_Update/ca
      -- 
    ca_11836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_2914_inst_ack_1, ack => cp_elements(826)); -- 
    -- CP-element group 827 transition  place  dead  bypass 
    -- predecessors 826 
    -- successors 45 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2922__entry__
      -- 	branch_block_stmt_1659/if_stmt_2916__exit__
      -- 	branch_block_stmt_1659/if_stmt_2916_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2916_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2916_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2922_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2922_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2922_dead_link/dead_transition
      -- 
    cp_elements(827) <= false;
    -- CP-element group 828 transition  output  bypass 
    -- predecessors 826 
    -- successors 829 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2916_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2916_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2916_eval_test/branch_req
      -- 
    cp_elements(828) <= cp_elements(826);
    branch_req_11844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => if_stmt_2916_branch_req_0); -- 
    -- CP-element group 829 branch  place  bypass 
    -- predecessors 828 
    -- successors 830 832 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_98_2917_place
      -- 
    cp_elements(829) <= cp_elements(828);
    -- CP-element group 830 transition  bypass 
    -- predecessors 829 
    -- successors 831 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2916_if_link/$entry
      -- 
    cp_elements(830) <= cp_elements(829);
    -- CP-element group 831 fork  transition  place  input  bypass 
    -- predecessors 830 
    -- successors 1900 1901 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2916_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2916_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_44_xx_xthread
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$entry
      -- 
    if_choice_transition_11849_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2916_branch_ack_1, ack => cp_elements(831)); -- 
    -- CP-element group 832 transition  bypass 
    -- predecessors 829 
    -- successors 833 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2916_else_link/$entry
      -- 
    cp_elements(832) <= cp_elements(829);
    -- CP-element group 833 transition  place  input  bypass 
    -- predecessors 832 
    -- successors 45 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2916_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2916_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_44_bb_45
      -- 	branch_block_stmt_1659/merge_stmt_2922_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_44_bb_45_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_44_bb_45_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2922_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2922_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2922_PhiAck/dummy
      -- 
    else_choice_transition_11853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2916_branch_ack_0, ack => cp_elements(833)); -- 
    -- CP-element group 834 fork  transition  bypass 
    -- predecessors 45 
    -- successors 835 836 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2928/$entry
      -- 
    cp_elements(834) <= cp_elements(45);
    -- CP-element group 835 transition  output  bypass 
    -- predecessors 834 
    -- successors 838 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Update/cr
      -- 
    cp_elements(835) <= cp_elements(834);
    cr_11875_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => SGT_f32_u1_2927_inst_req_1); -- 
    -- CP-element group 836 transition  output  bypass 
    -- predecessors 834 
    -- successors 837 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2928/R_iNsTr_97_2924_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2928/R_iNsTr_97_2924_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2928/R_iNsTr_97_2924_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2928/R_iNsTr_97_2924_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Sample/rr
      -- 
    cp_elements(836) <= cp_elements(834);
    rr_11870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(836), ack => SGT_f32_u1_2927_inst_req_0); -- 
    -- CP-element group 837 transition  input  bypass 
    -- predecessors 836 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Sample/ra
      -- 
    ra_11871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2927_inst_ack_0, ack => cp_elements(837)); -- 
    -- CP-element group 838 branch  transition  place  input  bypass 
    -- predecessors 835 
    -- successors 839 840 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2929__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2928__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2928/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2928/SGT_f32_u1_2927_Update/ca
      -- 
    ca_11876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f32_u1_2927_inst_ack_1, ack => cp_elements(838)); -- 
    -- CP-element group 839 transition  place  dead  bypass 
    -- predecessors 838 
    -- successors 46 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2935__entry__
      -- 	branch_block_stmt_1659/if_stmt_2929__exit__
      -- 	branch_block_stmt_1659/if_stmt_2929_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2929_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2929_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2935_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2935_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2935_dead_link/dead_transition
      -- 
    cp_elements(839) <= false;
    -- CP-element group 840 transition  output  bypass 
    -- predecessors 838 
    -- successors 841 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2929_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2929_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2929_eval_test/branch_req
      -- 
    cp_elements(840) <= cp_elements(838);
    branch_req_11884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => if_stmt_2929_branch_req_0); -- 
    -- CP-element group 841 branch  place  bypass 
    -- predecessors 840 
    -- successors 842 844 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_122_2930_place
      -- 
    cp_elements(841) <= cp_elements(840);
    -- CP-element group 842 transition  bypass 
    -- predecessors 841 
    -- successors 843 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2929_if_link/$entry
      -- 
    cp_elements(842) <= cp_elements(841);
    -- CP-element group 843 fork  transition  place  input  bypass 
    -- predecessors 842 
    -- successors 1903 1904 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2929_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2929_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_45_xx_xthread
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$entry
      -- 
    if_choice_transition_11889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2929_branch_ack_1, ack => cp_elements(843)); -- 
    -- CP-element group 844 transition  bypass 
    -- predecessors 841 
    -- successors 845 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2929_else_link/$entry
      -- 
    cp_elements(844) <= cp_elements(841);
    -- CP-element group 845 transition  place  input  bypass 
    -- predecessors 844 
    -- successors 46 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_2929_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2929_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_45_bb_46
      -- 	branch_block_stmt_1659/merge_stmt_2935_PhiReqMerge
      -- 	branch_block_stmt_1659/bb_45_bb_46_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_45_bb_46_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2935_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2935_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2935_PhiAck/dummy
      -- 
    else_choice_transition_11893_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2929_branch_ack_0, ack => cp_elements(845)); -- 
    -- CP-element group 846 fork  transition  bypass 
    -- predecessors 46 
    -- successors 847 848 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2941/$entry
      -- 
    cp_elements(846) <= cp_elements(46);
    -- CP-element group 847 transition  output  bypass 
    -- predecessors 846 
    -- successors 850 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Update/cr
      -- 
    cp_elements(847) <= cp_elements(846);
    cr_11915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(847), ack => EQ_f32_u1_2940_inst_req_1); -- 
    -- CP-element group 848 transition  output  bypass 
    -- predecessors 846 
    -- successors 849 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2941/R_iNsTr_97_2937_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2941/R_iNsTr_97_2937_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2941/R_iNsTr_97_2937_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2941/R_iNsTr_97_2937_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Sample/rr
      -- 
    cp_elements(848) <= cp_elements(846);
    rr_11910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => EQ_f32_u1_2940_inst_req_0); -- 
    -- CP-element group 849 transition  input  bypass 
    -- predecessors 848 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Sample/ra
      -- 
    ra_11911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2940_inst_ack_0, ack => cp_elements(849)); -- 
    -- CP-element group 850 branch  transition  place  input  bypass 
    -- predecessors 847 
    -- successors 851 852 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_2942__entry__
      -- 	branch_block_stmt_1659/assign_stmt_2941__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2941/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2941/EQ_f32_u1_2940_Update/ca
      -- 
    ca_11916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_f32_u1_2940_inst_ack_1, ack => cp_elements(850)); -- 
    -- CP-element group 851 transition  place  dead  bypass 
    -- predecessors 850 
    -- successors 47 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_2948__entry__
      -- 	branch_block_stmt_1659/if_stmt_2942__exit__
      -- 	branch_block_stmt_1659/if_stmt_2942_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_2942_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2942_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_2948_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_2948_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2948_dead_link/dead_transition
      -- 
    cp_elements(851) <= false;
    -- CP-element group 852 transition  output  bypass 
    -- predecessors 850 
    -- successors 853 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_2942_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_2942_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_2942_eval_test/branch_req
      -- 
    cp_elements(852) <= cp_elements(850);
    branch_req_11924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(852), ack => if_stmt_2942_branch_req_0); -- 
    -- CP-element group 853 branch  place  bypass 
    -- predecessors 852 
    -- successors 854 856 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_149_2943_place
      -- 
    cp_elements(853) <= cp_elements(852);
    -- CP-element group 854 transition  bypass 
    -- predecessors 853 
    -- successors 855 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2942_if_link/$entry
      -- 
    cp_elements(854) <= cp_elements(853);
    -- CP-element group 855 fork  transition  place  input  bypass 
    -- predecessors 854 
    -- successors 2159 2160 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2942_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2942_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/$entry
      -- 
    if_choice_transition_11929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2942_branch_ack_1, ack => cp_elements(855)); -- 
    -- CP-element group 856 transition  bypass 
    -- predecessors 853 
    -- successors 857 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_2942_else_link/$entry
      -- 
    cp_elements(856) <= cp_elements(853);
    -- CP-element group 857 fork  transition  place  input  bypass 
    -- predecessors 856 
    -- successors 1906 1908 
    -- members (8) 
      -- 	branch_block_stmt_1659/if_stmt_2942_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_2942_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/bb_46_xx_xthread
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$entry
      -- 
    else_choice_transition_11933_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2942_branch_ack_0, ack => cp_elements(857)); -- 
    -- CP-element group 858 fork  transition  bypass 
    -- predecessors 47 
    -- successors 859 860 863 866 869 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/$entry
      -- 
    cp_elements(858) <= cp_elements(47);
    -- CP-element group 859 transition  output  bypass 
    -- predecessors 858 
    -- successors 862 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_update_start_
      -- 
    cp_elements(859) <= cp_elements(858);
    cr_11955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(859), ack => type_cast_2962_inst_req_1); -- 
    -- CP-element group 860 transition  output  bypass 
    -- predecessors 858 
    -- successors 861 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35x_xin_2961_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35x_xin_2961_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35x_xin_2961_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35x_xin_2961_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_sample_start_
      -- 
    cp_elements(860) <= cp_elements(858);
    rr_11950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(860), ack => type_cast_2962_inst_req_0); -- 
    -- CP-element group 861 transition  input  bypass 
    -- predecessors 860 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_sample_completed_
      -- 
    ra_11951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2962_inst_ack_0, ack => cp_elements(861)); -- 
    -- CP-element group 862 transition  input  output  bypass 
    -- predecessors 859 
    -- successors 864 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35_2965_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35_2965_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35_2965_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/type_cast_2962_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_tmp10x_xi35_2965_sample_start_
      -- 
    ca_11956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2962_inst_ack_1, ack => cp_elements(862)); -- 
    rr_11968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(862), ack => SHL_u32_u32_2968_inst_req_0); -- 
    -- CP-element group 863 transition  output  bypass 
    -- predecessors 858 
    -- successors 865 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_update_start_
      -- 
    cp_elements(863) <= cp_elements(858);
    cr_11973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(863), ack => SHL_u32_u32_2968_inst_req_1); -- 
    -- CP-element group 864 transition  input  bypass 
    -- predecessors 862 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_sample_completed_
      -- 
    ra_11969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2968_inst_ack_0, ack => cp_elements(864)); -- 
    -- CP-element group 865 transition  input  output  bypass 
    -- predecessors 863 
    -- successors 867 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/SHL_u32_u32_2968_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_118_2971_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_118_2971_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_118_2971_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_118_2971_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Sample/rr
      -- 
    ca_11974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_2968_inst_ack_1, ack => cp_elements(865)); -- 
    rr_11986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(865), ack => AND_u32_u32_2974_inst_req_0); -- 
    -- CP-element group 866 transition  output  bypass 
    -- predecessors 858 
    -- successors 868 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Update/$entry
      -- 
    cp_elements(866) <= cp_elements(858);
    cr_11991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(866), ack => AND_u32_u32_2974_inst_req_1); -- 
    -- CP-element group 867 transition  input  bypass 
    -- predecessors 865 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Sample/ra
      -- 
    ra_11987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2974_inst_ack_0, ack => cp_elements(867)); -- 
    -- CP-element group 868 transition  input  output  bypass 
    -- predecessors 866 
    -- successors 870 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_119_2977_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_119_2977_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_119_2977_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/R_iNsTr_119_2977_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/AND_u32_u32_2974_Update/$exit
      -- 
    ca_11992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_2974_inst_ack_1, ack => cp_elements(868)); -- 
    rr_12004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => OR_u32_u32_2980_inst_req_0); -- 
    -- CP-element group 869 transition  output  bypass 
    -- predecessors 858 
    -- successors 871 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_update_start_
      -- 
    cp_elements(869) <= cp_elements(858);
    cr_12009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(869), ack => OR_u32_u32_2980_inst_req_1); -- 
    -- CP-element group 870 transition  input  bypass 
    -- predecessors 868 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Sample/$exit
      -- 
    ra_12005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2980_inst_ack_0, ack => cp_elements(870)); -- 
    -- CP-element group 871 transition  place  input  bypass 
    -- predecessors 869 
    -- successors 1934 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/OR_u32_u32_2980_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_2963_to_assign_stmt_2981/$exit
      -- 
    ca_12010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_2980_inst_ack_1, ack => cp_elements(871)); -- 
    -- CP-element group 872 fork  transition  bypass 
    -- predecessors 48 
    -- successors 873 874 877 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/$entry
      -- 
    cp_elements(872) <= cp_elements(48);
    -- CP-element group 873 transition  output  bypass 
    -- predecessors 872 
    -- successors 876 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Update/cr
      -- 
    cp_elements(873) <= cp_elements(872);
    cr_12030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(873), ack => LSHR_u32_u32_3002_inst_req_1); -- 
    -- CP-element group 874 transition  output  bypass 
    -- predecessors 872 
    -- successors 875 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_xx_x016x_xix_xi_2999_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_xx_x016x_xix_xi_2999_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_xx_x016x_xix_xi_2999_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_xx_x016x_xix_xi_2999_update_start_
      -- 
    cp_elements(874) <= cp_elements(872);
    rr_12025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => LSHR_u32_u32_3002_inst_req_0); -- 
    -- CP-element group 875 transition  input  bypass 
    -- predecessors 874 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_sample_completed_
      -- 
    ra_12026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3002_inst_ack_0, ack => cp_elements(875)); -- 
    -- CP-element group 876 transition  input  output  bypass 
    -- predecessors 873 
    -- successors 878 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/LSHR_u32_u32_3002_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_iNsTr_146_3005_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_iNsTr_146_3005_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_iNsTr_146_3005_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/R_iNsTr_146_3005_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Sample/rr
      -- 
    ca_12031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3002_inst_ack_1, ack => cp_elements(876)); -- 
    rr_12043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(876), ack => UGT_u32_u1_3008_inst_req_0); -- 
    -- CP-element group 877 transition  output  bypass 
    -- predecessors 872 
    -- successors 879 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Update/cr
      -- 
    cp_elements(877) <= cp_elements(872);
    cr_12048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(877), ack => UGT_u32_u1_3008_inst_req_1); -- 
    -- CP-element group 878 transition  input  bypass 
    -- predecessors 876 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Sample/ra
      -- 
    ra_12044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3008_inst_ack_0, ack => cp_elements(878)); -- 
    -- CP-element group 879 branch  transition  place  input  bypass 
    -- predecessors 877 
    -- successors 880 881 
    -- members (6) 
      -- 	branch_block_stmt_1659/if_stmt_3010__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3003_to_assign_stmt_3009/UGT_u32_u1_3008_Update/ca
      -- 
    ca_12049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u32_u1_3008_inst_ack_1, ack => cp_elements(879)); -- 
    -- CP-element group 880 transition  place  dead  bypass 
    -- predecessors 879 
    -- successors 49 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3016__entry__
      -- 	branch_block_stmt_1659/if_stmt_3010__exit__
      -- 	branch_block_stmt_1659/if_stmt_3010_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_3010_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3010_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_3016_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3016_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3016_dead_link/dead_transition
      -- 
    cp_elements(880) <= false;
    -- CP-element group 881 transition  output  bypass 
    -- predecessors 879 
    -- successors 882 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3010_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_3010_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_3010_eval_test/branch_req
      -- 
    cp_elements(881) <= cp_elements(879);
    branch_req_12057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(881), ack => if_stmt_3010_branch_req_0); -- 
    -- CP-element group 882 branch  place  bypass 
    -- predecessors 881 
    -- successors 883 885 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_147_3011_place
      -- 
    cp_elements(882) <= cp_elements(881);
    -- CP-element group 883 transition  bypass 
    -- predecessors 882 
    -- successors 884 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3010_if_link/$entry
      -- 
    cp_elements(883) <= cp_elements(882);
    -- CP-element group 884 transition  place  input  bypass 
    -- predecessors 883 
    -- successors 49 
    -- members (9) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader
      -- 	branch_block_stmt_1659/if_stmt_3010_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3010_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/merge_stmt_3016_PhiReqMerge
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_bbx_xnphx_xix_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3016_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3016_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3016_PhiAck/dummy
      -- 
    if_choice_transition_12062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3010_branch_ack_1, ack => cp_elements(884)); -- 
    -- CP-element group 885 transition  bypass 
    -- predecessors 882 
    -- successors 886 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3010_else_link/$entry
      -- 
    cp_elements(885) <= cp_elements(882);
    -- CP-element group 886 transition  place  input  bypass 
    -- predecessors 885 
    -- successors 2005 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_3010_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3010_else_link/else_choice_transition
      -- 
    else_choice_transition_12066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3010_branch_ack_0, ack => cp_elements(886)); -- 
    -- CP-element group 887 fork  transition  bypass 
    -- predecessors 50 
    -- successors 888 889 892 893 897 898 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/$entry
      -- 
    cp_elements(887) <= cp_elements(50);
    -- CP-element group 888 transition  output  bypass 
    -- predecessors 887 
    -- successors 891 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Update/cr
      -- 
    cp_elements(888) <= cp_elements(887);
    cr_12088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(888), ack => SHL_u32_u32_3038_inst_req_1); -- 
    -- CP-element group 889 transition  output  bypass 
    -- predecessors 887 
    -- successors 890 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_shifted_divisorx_x03x_xix_xi_3035_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_shifted_divisorx_x03x_xix_xi_3035_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_shifted_divisorx_x03x_xix_xi_3035_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_shifted_divisorx_x03x_xix_xi_3035_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Sample/rr
      -- 
    cp_elements(889) <= cp_elements(887);
    rr_12083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(889), ack => SHL_u32_u32_3038_inst_req_0); -- 
    -- CP-element group 890 transition  input  bypass 
    -- predecessors 889 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Sample/ra
      -- 
    ra_12084_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3038_inst_ack_0, ack => cp_elements(890)); -- 
    -- CP-element group 891 transition  input  bypass 
    -- predecessors 888 
    -- successors 896 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3038_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_190_3047_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_190_3047_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_190_3047_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_190_3047_update_completed_
      -- 
    ca_12089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3038_inst_ack_1, ack => cp_elements(891)); -- 
    -- CP-element group 892 transition  output  bypass 
    -- predecessors 887 
    -- successors 895 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Update/cr
      -- 
    cp_elements(892) <= cp_elements(887);
    cr_12106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(892), ack => SHL_u32_u32_3044_inst_req_1); -- 
    -- CP-element group 893 transition  output  bypass 
    -- predecessors 887 
    -- successors 894 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_curr_quotientx_x02x_xix_xi_3041_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_curr_quotientx_x02x_xix_xi_3041_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_curr_quotientx_x02x_xix_xi_3041_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_curr_quotientx_x02x_xix_xi_3041_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Sample/rr
      -- 
    cp_elements(893) <= cp_elements(887);
    rr_12101_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(893), ack => SHL_u32_u32_3044_inst_req_0); -- 
    -- CP-element group 894 transition  input  bypass 
    -- predecessors 893 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Sample/ra
      -- 
    ra_12102_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3044_inst_ack_0, ack => cp_elements(894)); -- 
    -- CP-element group 895 transition  input  bypass 
    -- predecessors 892 
    -- successors 901 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/SHL_u32_u32_3044_Update/ca
      -- 
    ca_12107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3044_inst_ack_1, ack => cp_elements(895)); -- 
    -- CP-element group 896 join  transition  output  bypass 
    -- predecessors 891 898 
    -- successors 899 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Sample/rr
      -- 
    cp_element_group_896: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_896"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(891) & cp_elements(898);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(896), clk => clk, reset => reset); --
    end block;
    rr_12123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(896), ack => ULT_u32_u1_3049_inst_req_0); -- 
    -- CP-element group 897 transition  output  bypass 
    -- predecessors 887 
    -- successors 900 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Update/cr
      -- 
    cp_elements(897) <= cp_elements(887);
    cr_12128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(897), ack => ULT_u32_u1_3049_inst_req_1); -- 
    -- CP-element group 898 transition  bypass 
    -- predecessors 887 
    -- successors 896 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_146_3048_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_146_3048_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_146_3048_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/R_iNsTr_146_3048_update_completed_
      -- 
    cp_elements(898) <= cp_elements(887);
    -- CP-element group 899 transition  input  bypass 
    -- predecessors 896 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Sample/ra
      -- 
    ra_12124_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3049_inst_ack_0, ack => cp_elements(899)); -- 
    -- CP-element group 900 transition  input  bypass 
    -- predecessors 897 
    -- successors 901 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/ULT_u32_u1_3049_Update/ca
      -- 
    ca_12129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3049_inst_ack_1, ack => cp_elements(900)); -- 
    -- CP-element group 901 join  transition  bypass 
    -- predecessors 895 900 
    -- successors 51 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3039_to_assign_stmt_3050/$exit
      -- 
    cp_element_group_901: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_901"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(895) & cp_elements(900);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(901), clk => clk, reset => reset); --
    end block;
    -- CP-element group 902 transition  place  dead  bypass 
    -- predecessors 51 
    -- successors 52 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3057__entry__
      -- 	branch_block_stmt_1659/if_stmt_3051__exit__
      -- 	branch_block_stmt_1659/if_stmt_3051_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_3051_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3051_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_3057_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3057_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3057_dead_link/dead_transition
      -- 
    cp_elements(902) <= false;
    -- CP-element group 903 transition  output  bypass 
    -- predecessors 51 
    -- successors 904 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3051_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_3051_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_3051_eval_test/branch_req
      -- 
    cp_elements(903) <= cp_elements(51);
    branch_req_12137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(903), ack => if_stmt_3051_branch_req_0); -- 
    -- CP-element group 904 branch  place  bypass 
    -- predecessors 903 
    -- successors 905 907 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_192_3052_place
      -- 
    cp_elements(904) <= cp_elements(903);
    -- CP-element group 905 transition  bypass 
    -- predecessors 904 
    -- successors 906 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3051_if_link/$entry
      -- 
    cp_elements(905) <= cp_elements(904);
    -- CP-element group 906 transition  place  input  bypass 
    -- predecessors 905 
    -- successors 1957 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_3051_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3051_if_link/if_choice_transition
      -- 
    if_choice_transition_12142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3051_branch_ack_1, ack => cp_elements(906)); -- 
    -- CP-element group 907 transition  bypass 
    -- predecessors 904 
    -- successors 908 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3051_else_link/$entry
      -- 
    cp_elements(907) <= cp_elements(904);
    -- CP-element group 908 transition  place  input  bypass 
    -- predecessors 907 
    -- successors 1986 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit
      -- 	branch_block_stmt_1659/if_stmt_3051_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3051_else_link/else_choice_transition
      -- 
    else_choice_transition_12146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3051_branch_ack_0, ack => cp_elements(908)); -- 
    -- CP-element group 909 fork  transition  bypass 
    -- predecessors 53 
    -- successors 911 912 913 917 918 919 922 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/$entry
      -- 
    cp_elements(909) <= cp_elements(53);
    -- CP-element group 910 join  transition  output  bypass 
    -- predecessors 912 913 
    -- successors 914 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Sample/rr
      -- 
    cp_element_group_910: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_910"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(912) & cp_elements(913);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(910), clk => clk, reset => reset); --
    end block;
    rr_12167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(910), ack => ADD_u32_u32_3087_inst_req_0); -- 
    -- CP-element group 911 transition  output  bypass 
    -- predecessors 909 
    -- successors 915 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Update/cr
      -- 
    cp_elements(911) <= cp_elements(909);
    cr_12172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => ADD_u32_u32_3087_inst_req_1); -- 
    -- CP-element group 912 transition  bypass 
    -- predecessors 909 
    -- successors 910 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_curr_quotientx_x0x_xlcssax_xix_xi_3085_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_curr_quotientx_x0x_xlcssax_xix_xi_3085_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_curr_quotientx_x0x_xlcssax_xix_xi_3085_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_curr_quotientx_x0x_xlcssax_xix_xi_3085_update_completed_
      -- 
    cp_elements(912) <= cp_elements(909);
    -- CP-element group 913 transition  bypass 
    -- predecessors 909 
    -- successors 910 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_quotientx_x05x_xix_xi_3086_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_quotientx_x05x_xix_xi_3086_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_quotientx_x05x_xix_xi_3086_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_quotientx_x05x_xix_xi_3086_update_completed_
      -- 
    cp_elements(913) <= cp_elements(909);
    -- CP-element group 914 transition  input  bypass 
    -- predecessors 910 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Sample/ra
      -- 
    ra_12168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3087_inst_ack_0, ack => cp_elements(914)); -- 
    -- CP-element group 915 transition  input  bypass 
    -- predecessors 911 
    -- successors 925 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ADD_u32_u32_3087_Update/ca
      -- 
    ca_12173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3087_inst_ack_1, ack => cp_elements(915)); -- 
    -- CP-element group 916 join  transition  output  bypass 
    -- predecessors 918 919 
    -- successors 920 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Sample/rr
      -- 
    cp_element_group_916: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_916"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(918) & cp_elements(919);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(916), clk => clk, reset => reset); --
    end block;
    rr_12189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(916), ack => SUB_u32_u32_3092_inst_req_0); -- 
    -- CP-element group 917 transition  output  bypass 
    -- predecessors 909 
    -- successors 921 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Update/cr
      -- 
    cp_elements(917) <= cp_elements(909);
    cr_12194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(917), ack => SUB_u32_u32_3092_inst_req_1); -- 
    -- CP-element group 918 transition  bypass 
    -- predecessors 909 
    -- successors 916 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_xx_x016x_xix_xi_3090_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_xx_x016x_xix_xi_3090_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_xx_x016x_xix_xi_3090_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_xx_x016x_xix_xi_3090_update_completed_
      -- 
    cp_elements(918) <= cp_elements(909);
    -- CP-element group 919 transition  bypass 
    -- predecessors 909 
    -- successors 916 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_shifted_divisorx_x0x_xlcssax_xix_xi_3091_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_shifted_divisorx_x0x_xlcssax_xix_xi_3091_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_shifted_divisorx_x0x_xlcssax_xix_xi_3091_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_shifted_divisorx_x0x_xlcssax_xix_xi_3091_update_completed_
      -- 
    cp_elements(919) <= cp_elements(909);
    -- CP-element group 920 transition  input  bypass 
    -- predecessors 916 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Sample/ra
      -- 
    ra_12190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3092_inst_ack_0, ack => cp_elements(920)); -- 
    -- CP-element group 921 transition  input  output  bypass 
    -- predecessors 917 
    -- successors 923 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/SUB_u32_u32_3092_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_iNsTr_170_3095_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_iNsTr_170_3095_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_iNsTr_170_3095_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/R_iNsTr_170_3095_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Sample/rr
      -- 
    ca_12195_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3092_inst_ack_1, ack => cp_elements(921)); -- 
    rr_12207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(921), ack => ULT_u32_u1_3098_inst_req_0); -- 
    -- CP-element group 922 transition  output  bypass 
    -- predecessors 909 
    -- successors 924 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Update/cr
      -- 
    cp_elements(922) <= cp_elements(909);
    cr_12212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(922), ack => ULT_u32_u1_3098_inst_req_1); -- 
    -- CP-element group 923 transition  input  bypass 
    -- predecessors 921 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Sample/ra
      -- 
    ra_12208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3098_inst_ack_0, ack => cp_elements(923)); -- 
    -- CP-element group 924 transition  input  bypass 
    -- predecessors 922 
    -- successors 925 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/ULT_u32_u1_3098_Update/ca
      -- 
    ca_12213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_3098_inst_ack_1, ack => cp_elements(924)); -- 
    -- CP-element group 925 join  transition  bypass 
    -- predecessors 915 924 
    -- successors 54 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3088_to_assign_stmt_3099/$exit
      -- 
    cp_element_group_925: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_925"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(915) & cp_elements(924);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 926 transition  place  dead  bypass 
    -- predecessors 54 
    -- successors 55 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3106__entry__
      -- 	branch_block_stmt_1659/if_stmt_3100__exit__
      -- 	branch_block_stmt_1659/if_stmt_3100_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_3100_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3100_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_3106_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3106_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3106_dead_link/dead_transition
      -- 
    cp_elements(926) <= false;
    -- CP-element group 927 transition  output  bypass 
    -- predecessors 54 
    -- successors 928 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3100_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_3100_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_3100_eval_test/branch_req
      -- 
    cp_elements(927) <= cp_elements(54);
    branch_req_12221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(927), ack => if_stmt_3100_branch_req_0); -- 
    -- CP-element group 928 branch  place  bypass 
    -- predecessors 927 
    -- successors 929 931 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_iNsTr_171_3101_place
      -- 
    cp_elements(928) <= cp_elements(927);
    -- CP-element group 929 transition  bypass 
    -- predecessors 928 
    -- successors 930 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3100_if_link/$entry
      -- 
    cp_elements(929) <= cp_elements(928);
    -- CP-element group 930 fork  transition  place  input  bypass 
    -- predecessors 929 
    -- successors 2034 2036 
    -- members (8) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi
      -- 	branch_block_stmt_1659/if_stmt_3100_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3100_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/$entry
      -- 
    if_choice_transition_12226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3100_branch_ack_1, ack => cp_elements(930)); -- 
    -- CP-element group 931 transition  bypass 
    -- predecessors 928 
    -- successors 932 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3100_else_link/$entry
      -- 
    cp_elements(931) <= cp_elements(928);
    -- CP-element group 932 transition  place  input  bypass 
    -- predecessors 931 
    -- successors 1914 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi
      -- 	branch_block_stmt_1659/if_stmt_3100_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3100_else_link/else_choice_transition
      -- 
    else_choice_transition_12230_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3100_branch_ack_0, ack => cp_elements(932)); -- 
    -- CP-element group 933 fork  transition  bypass 
    -- predecessors 55 
    -- successors 934 935 938 939 942 945 948 949 952 955 956 962 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/$entry
      -- 
    cp_elements(933) <= cp_elements(55);
    -- CP-element group 934 transition  output  bypass 
    -- predecessors 933 
    -- successors 937 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Update/cr
      -- 
    cp_elements(934) <= cp_elements(933);
    cr_12252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(934), ack => LSHR_u32_u32_3116_inst_req_1); -- 
    -- CP-element group 935 transition  output  bypass 
    -- predecessors 933 
    -- successors 936 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3113_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3113_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3113_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3113_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Sample/rr
      -- 
    cp_elements(935) <= cp_elements(933);
    rr_12247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => LSHR_u32_u32_3116_inst_req_0); -- 
    -- CP-element group 936 transition  input  bypass 
    -- predecessors 935 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Sample/ra
      -- 
    ra_12248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3116_inst_ack_0, ack => cp_elements(936)); -- 
    -- CP-element group 937 transition  input  output  bypass 
    -- predecessors 934 
    -- successors 943 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/LSHR_u32_u32_3116_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_194_3125_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_194_3125_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_194_3125_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_194_3125_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Sample/rr
      -- 
    ca_12253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_3116_inst_ack_1, ack => cp_elements(937)); -- 
    rr_12283_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(937), ack => AND_u32_u32_3128_inst_req_0); -- 
    -- CP-element group 938 transition  output  bypass 
    -- predecessors 933 
    -- successors 941 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Update/cr
      -- 
    cp_elements(938) <= cp_elements(933);
    cr_12270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(938), ack => AND_u32_u32_3122_inst_req_1); -- 
    -- CP-element group 939 transition  output  bypass 
    -- predecessors 933 
    -- successors 940 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3119_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3119_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3119_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_tmp10x_xi35_3119_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Sample/rr
      -- 
    cp_elements(939) <= cp_elements(933);
    rr_12265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => AND_u32_u32_3122_inst_req_0); -- 
    -- CP-element group 940 transition  input  bypass 
    -- predecessors 939 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Sample/ra
      -- 
    ra_12266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3122_inst_ack_0, ack => cp_elements(940)); -- 
    -- CP-element group 941 transition  input  bypass 
    -- predecessors 938 
    -- successors 965 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3122_Update/ca
      -- 
    ca_12271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3122_inst_ack_1, ack => cp_elements(941)); -- 
    -- CP-element group 942 transition  output  bypass 
    -- predecessors 933 
    -- successors 944 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Update/cr
      -- 
    cp_elements(942) <= cp_elements(933);
    cr_12288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(942), ack => AND_u32_u32_3128_inst_req_1); -- 
    -- CP-element group 943 transition  input  bypass 
    -- predecessors 937 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Sample/ra
      -- 
    ra_12284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3128_inst_ack_0, ack => cp_elements(943)); -- 
    -- CP-element group 944 transition  input  output  bypass 
    -- predecessors 942 
    -- successors 946 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3128_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_196_3131_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_196_3131_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_196_3131_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_196_3131_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Sample/rr
      -- 
    ca_12289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3128_inst_ack_1, ack => cp_elements(944)); -- 
    rr_12301_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => ADD_u32_u32_3134_inst_req_0); -- 
    -- CP-element group 945 transition  output  bypass 
    -- predecessors 933 
    -- successors 947 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Update/cr
      -- 
    cp_elements(945) <= cp_elements(933);
    cr_12306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(945), ack => ADD_u32_u32_3134_inst_req_1); -- 
    -- CP-element group 946 transition  input  bypass 
    -- predecessors 944 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Sample/ra
      -- 
    ra_12302_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3134_inst_ack_0, ack => cp_elements(946)); -- 
    -- CP-element group 947 transition  input  bypass 
    -- predecessors 945 
    -- successors 965 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/ADD_u32_u32_3134_Update/ca
      -- 
    ca_12307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3134_inst_ack_1, ack => cp_elements(947)); -- 
    -- CP-element group 948 transition  output  bypass 
    -- predecessors 933 
    -- successors 951 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Update/cr
      -- 
    cp_elements(948) <= cp_elements(933);
    cr_12324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(948), ack => AND_u32_u32_3140_inst_req_1); -- 
    -- CP-element group 949 transition  output  bypass 
    -- predecessors 933 
    -- successors 950 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3137_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3137_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3137_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3137_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Sample/rr
      -- 
    cp_elements(949) <= cp_elements(933);
    rr_12319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => AND_u32_u32_3140_inst_req_0); -- 
    -- CP-element group 950 transition  input  bypass 
    -- predecessors 949 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Sample/ra
      -- 
    ra_12320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3140_inst_ack_0, ack => cp_elements(950)); -- 
    -- CP-element group 951 transition  input  output  bypass 
    -- predecessors 948 
    -- successors 953 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u32_u32_3140_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_198_3143_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_198_3143_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_198_3143_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_198_3143_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Sample/rr
      -- 
    ca_12325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3140_inst_ack_1, ack => cp_elements(951)); -- 
    rr_12337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(951), ack => EQ_u32_u1_3146_inst_req_0); -- 
    -- CP-element group 952 transition  output  bypass 
    -- predecessors 933 
    -- successors 954 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Update/cr
      -- 
    cp_elements(952) <= cp_elements(933);
    cr_12342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(952), ack => EQ_u32_u1_3146_inst_req_1); -- 
    -- CP-element group 953 transition  input  bypass 
    -- predecessors 951 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Sample/ra
      -- 
    ra_12338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3146_inst_ack_0, ack => cp_elements(953)); -- 
    -- CP-element group 954 transition  input  bypass 
    -- predecessors 952 
    -- successors 961 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/EQ_u32_u1_3146_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_199_3157_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_199_3157_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_199_3157_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_199_3157_update_completed_
      -- 
    ca_12343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3146_inst_ack_1, ack => cp_elements(954)); -- 
    -- CP-element group 955 transition  output  bypass 
    -- predecessors 933 
    -- successors 960 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Update/cr
      -- 
    cp_elements(955) <= cp_elements(933);
    cr_12374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => NEQ_i32_u1_3154_inst_req_1); -- 
    -- CP-element group 956 transition  output  bypass 
    -- predecessors 933 
    -- successors 957 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3149_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3149_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3149_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_xx_xlcssa4_3149_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Sample/rr
      -- 
    cp_elements(956) <= cp_elements(933);
    rr_12359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(956), ack => type_cast_3150_inst_req_0); -- 
    -- CP-element group 957 transition  input  output  bypass 
    -- predecessors 956 
    -- successors 958 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Update/cr
      -- 
    ra_12360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3150_inst_ack_0, ack => cp_elements(957)); -- 
    cr_12364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(957), ack => type_cast_3150_inst_req_1); -- 
    -- CP-element group 958 transition  input  output  bypass 
    -- predecessors 957 
    -- successors 959 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/type_cast_3150_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Sample/rr
      -- 
    ca_12365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3150_inst_ack_1, ack => cp_elements(958)); -- 
    rr_12369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(958), ack => NEQ_i32_u1_3154_inst_req_0); -- 
    -- CP-element group 959 transition  input  bypass 
    -- predecessors 958 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Sample/ra
      -- 
    ra_12370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3154_inst_ack_0, ack => cp_elements(959)); -- 
    -- CP-element group 960 transition  input  bypass 
    -- predecessors 955 
    -- successors 961 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/NEQ_i32_u1_3154_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_200_3158_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_200_3158_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_200_3158_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/R_iNsTr_200_3158_update_completed_
      -- 
    ca_12375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3154_inst_ack_1, ack => cp_elements(960)); -- 
    -- CP-element group 961 join  transition  output  bypass 
    -- predecessors 954 960 
    -- successors 963 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Sample/rr
      -- 
    cp_element_group_961: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_961"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(954) & cp_elements(960);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(961), clk => clk, reset => reset); --
    end block;
    rr_12391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => AND_u1_u1_3159_inst_req_0); -- 
    -- CP-element group 962 transition  output  bypass 
    -- predecessors 933 
    -- successors 964 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Update/cr
      -- 
    cp_elements(962) <= cp_elements(933);
    cr_12396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => AND_u1_u1_3159_inst_req_1); -- 
    -- CP-element group 963 transition  input  bypass 
    -- predecessors 961 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Sample/ra
      -- 
    ra_12392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3159_inst_ack_0, ack => cp_elements(963)); -- 
    -- CP-element group 964 transition  input  bypass 
    -- predecessors 962 
    -- successors 965 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/AND_u1_u1_3159_Update/ca
      -- 
    ca_12397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3159_inst_ack_1, ack => cp_elements(964)); -- 
    -- CP-element group 965 join  transition  bypass 
    -- predecessors 941 947 964 
    -- successors 56 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3117_to_assign_stmt_3160/$exit
      -- 
    cp_element_group_965: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_965"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(941) & cp_elements(947) & cp_elements(964);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(965), clk => clk, reset => reset); --
    end block;
    -- CP-element group 966 transition  place  dead  bypass 
    -- predecessors 56 
    -- successors 57 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3167__entry__
      -- 	branch_block_stmt_1659/if_stmt_3161__exit__
      -- 	branch_block_stmt_1659/if_stmt_3161_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_3161_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3161_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_3167_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3167_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3167_dead_link/dead_transition
      -- 
    cp_elements(966) <= false;
    -- CP-element group 967 transition  output  bypass 
    -- predecessors 56 
    -- successors 968 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3161_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_3161_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_3161_eval_test/branch_req
      -- 
    cp_elements(967) <= cp_elements(56);
    branch_req_12405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(967), ack => if_stmt_3161_branch_req_0); -- 
    -- CP-element group 968 branch  place  bypass 
    -- predecessors 967 
    -- successors 969 971 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcond11x_xi_3162_place
      -- 
    cp_elements(968) <= cp_elements(967);
    -- CP-element group 969 transition  bypass 
    -- predecessors 968 
    -- successors 970 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3161_if_link/$entry
      -- 
    cp_elements(969) <= cp_elements(968);
    -- CP-element group 970 transition  place  input  bypass 
    -- predecessors 969 
    -- successors 57 
    -- members (9) 
      -- 	branch_block_stmt_1659/if_stmt_3161_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3161_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader
      -- 	branch_block_stmt_1659/merge_stmt_3167_PhiReqMerge
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_udiv32x_xexitx_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3167_PhiAck/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3167_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3167_PhiAck/dummy
      -- 
    if_choice_transition_12410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3161_branch_ack_1, ack => cp_elements(970)); -- 
    -- CP-element group 971 transition  bypass 
    -- predecessors 968 
    -- successors 972 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3161_else_link/$entry
      -- 
    cp_elements(971) <= cp_elements(968);
    -- CP-element group 972 transition  place  input  bypass 
    -- predecessors 971 
    -- successors 2102 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3161_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3161_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi
      -- 
    else_choice_transition_12414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3161_branch_ack_0, ack => cp_elements(972)); -- 
    -- CP-element group 973 fork  transition  bypass 
    -- predecessors 58 
    -- successors 974 975 978 982 985 992 995 996 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/$entry
      -- 
    cp_elements(973) <= cp_elements(58);
    -- CP-element group 974 transition  output  bypass 
    -- predecessors 973 
    -- successors 977 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Update/cr
      -- 
    cp_elements(974) <= cp_elements(973);
    cr_12436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(974), ack => SHL_u32_u32_3188_inst_req_1); -- 
    -- CP-element group 975 transition  output  bypass 
    -- predecessors 973 
    -- successors 976 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_tempx_x012x_xi_3185_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_tempx_x012x_xi_3185_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_tempx_x012x_xi_3185_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_tempx_x012x_xi_3185_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Sample/rr
      -- 
    cp_elements(975) <= cp_elements(973);
    rr_12431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(975), ack => SHL_u32_u32_3188_inst_req_0); -- 
    -- CP-element group 976 transition  input  bypass 
    -- predecessors 975 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Sample/ra
      -- 
    ra_12432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3188_inst_ack_0, ack => cp_elements(976)); -- 
    -- CP-element group 977 fork  transition  input  bypass 
    -- predecessors 974 
    -- successors 979 986 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/SHL_u32_u32_3188_Update/ca
      -- 
    ca_12437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3188_inst_ack_1, ack => cp_elements(977)); -- 
    -- CP-element group 978 transition  output  bypass 
    -- predecessors 973 
    -- successors 981 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Update/cr
      -- 
    cp_elements(978) <= cp_elements(973);
    cr_12454_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(978), ack => AND_u32_u32_3194_inst_req_1); -- 
    -- CP-element group 979 transition  output  bypass 
    -- predecessors 977 
    -- successors 980 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3191_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3191_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3191_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3191_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Sample/rr
      -- 
    cp_elements(979) <= cp_elements(977);
    rr_12449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(979), ack => AND_u32_u32_3194_inst_req_0); -- 
    -- CP-element group 980 transition  input  bypass 
    -- predecessors 979 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Sample/ra
      -- 
    ra_12450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3194_inst_ack_0, ack => cp_elements(980)); -- 
    -- CP-element group 981 transition  input  output  bypass 
    -- predecessors 978 
    -- successors 983 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u32_u32_3194_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_213_3197_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_213_3197_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_213_3197_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_213_3197_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Sample/rr
      -- 
    ca_12455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3194_inst_ack_1, ack => cp_elements(981)); -- 
    rr_12467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(981), ack => EQ_u32_u1_3200_inst_req_0); -- 
    -- CP-element group 982 transition  output  bypass 
    -- predecessors 973 
    -- successors 984 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Update/cr
      -- 
    cp_elements(982) <= cp_elements(973);
    cr_12472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(982), ack => EQ_u32_u1_3200_inst_req_1); -- 
    -- CP-element group 983 transition  input  bypass 
    -- predecessors 981 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Sample/ra
      -- 
    ra_12468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3200_inst_ack_0, ack => cp_elements(983)); -- 
    -- CP-element group 984 transition  input  bypass 
    -- predecessors 982 
    -- successors 991 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/EQ_u32_u1_3200_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_214_3211_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_214_3211_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_214_3211_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_214_3211_update_completed_
      -- 
    ca_12473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_3200_inst_ack_1, ack => cp_elements(984)); -- 
    -- CP-element group 985 transition  output  bypass 
    -- predecessors 973 
    -- successors 990 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Update/cr
      -- 
    cp_elements(985) <= cp_elements(973);
    cr_12504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(985), ack => NEQ_i32_u1_3208_inst_req_1); -- 
    -- CP-element group 986 transition  output  bypass 
    -- predecessors 977 
    -- successors 987 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3203_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3203_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3203_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_212_3203_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Sample/rr
      -- 
    cp_elements(986) <= cp_elements(977);
    rr_12489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(986), ack => type_cast_3204_inst_req_0); -- 
    -- CP-element group 987 transition  input  output  bypass 
    -- predecessors 986 
    -- successors 988 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Update/cr
      -- 
    ra_12490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3204_inst_ack_0, ack => cp_elements(987)); -- 
    cr_12494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(987), ack => type_cast_3204_inst_req_1); -- 
    -- CP-element group 988 transition  input  output  bypass 
    -- predecessors 987 
    -- successors 989 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/type_cast_3204_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Sample/rr
      -- 
    ca_12495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3204_inst_ack_1, ack => cp_elements(988)); -- 
    rr_12499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(988), ack => NEQ_i32_u1_3208_inst_req_0); -- 
    -- CP-element group 989 transition  input  bypass 
    -- predecessors 988 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Sample/ra
      -- 
    ra_12500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3208_inst_ack_0, ack => cp_elements(989)); -- 
    -- CP-element group 990 transition  input  bypass 
    -- predecessors 985 
    -- successors 991 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/NEQ_i32_u1_3208_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_215_3212_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_215_3212_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_215_3212_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_215_3212_update_completed_
      -- 
    ca_12505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => NEQ_i32_u1_3208_inst_ack_1, ack => cp_elements(990)); -- 
    -- CP-element group 991 join  transition  output  bypass 
    -- predecessors 984 990 
    -- successors 993 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Sample/rr
      -- 
    cp_element_group_991: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_991"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(984) & cp_elements(990);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(991), clk => clk, reset => reset); --
    end block;
    rr_12521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(991), ack => AND_u1_u1_3213_inst_req_0); -- 
    -- CP-element group 992 transition  output  bypass 
    -- predecessors 973 
    -- successors 994 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Update/cr
      -- 
    cp_elements(992) <= cp_elements(973);
    cr_12526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(992), ack => AND_u1_u1_3213_inst_req_1); -- 
    -- CP-element group 993 transition  input  bypass 
    -- predecessors 991 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Sample/ra
      -- 
    ra_12522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3213_inst_ack_0, ack => cp_elements(993)); -- 
    -- CP-element group 994 transition  input  bypass 
    -- predecessors 992 
    -- successors 999 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/AND_u1_u1_3213_Update/ca
      -- 
    ca_12527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3213_inst_ack_1, ack => cp_elements(994)); -- 
    -- CP-element group 995 transition  output  bypass 
    -- predecessors 973 
    -- successors 998 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Update/cr
      -- 
    cp_elements(995) <= cp_elements(973);
    cr_12544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(995), ack => ADD_u32_u32_3219_inst_req_1); -- 
    -- CP-element group 996 transition  output  bypass 
    -- predecessors 973 
    -- successors 997 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_211_3216_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_211_3216_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_211_3216_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/R_iNsTr_211_3216_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Sample/rr
      -- 
    cp_elements(996) <= cp_elements(973);
    rr_12539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(996), ack => ADD_u32_u32_3219_inst_req_0); -- 
    -- CP-element group 997 transition  input  bypass 
    -- predecessors 996 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Sample/ra
      -- 
    ra_12540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3219_inst_ack_0, ack => cp_elements(997)); -- 
    -- CP-element group 998 transition  input  bypass 
    -- predecessors 995 
    -- successors 999 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/ADD_u32_u32_3219_Update/ca
      -- 
    ca_12545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3219_inst_ack_1, ack => cp_elements(998)); -- 
    -- CP-element group 999 join  transition  bypass 
    -- predecessors 994 998 
    -- successors 59 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3189_to_assign_stmt_3220/$exit
      -- 
    cp_element_group_999: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 20) := "cp_element_group_999"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(994) & cp_elements(998);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(999), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1000 transition  place  dead  bypass 
    -- predecessors 59 
    -- successors 60 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3227__entry__
      -- 	branch_block_stmt_1659/if_stmt_3221__exit__
      -- 	branch_block_stmt_1659/if_stmt_3221_dead_link/$entry
      -- 	branch_block_stmt_1659/if_stmt_3221_dead_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3221_dead_link/dead_transition
      -- 	branch_block_stmt_1659/merge_stmt_3227_dead_link/$entry
      -- 	branch_block_stmt_1659/merge_stmt_3227_dead_link/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3227_dead_link/dead_transition
      -- 
    cp_elements(1000) <= false;
    -- CP-element group 1001 transition  output  bypass 
    -- predecessors 59 
    -- successors 1002 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3221_eval_test/$entry
      -- 	branch_block_stmt_1659/if_stmt_3221_eval_test/$exit
      -- 	branch_block_stmt_1659/if_stmt_3221_eval_test/branch_req
      -- 
    cp_elements(1001) <= cp_elements(59);
    branch_req_12553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1001), ack => if_stmt_3221_branch_req_0); -- 
    -- CP-element group 1002 branch  place  bypass 
    -- predecessors 1001 
    -- successors 1003 1005 
    -- members (1) 
      -- 	branch_block_stmt_1659/R_orx_xcondx_xi_3222_place
      -- 
    cp_elements(1002) <= cp_elements(1001);
    -- CP-element group 1003 transition  bypass 
    -- predecessors 1002 
    -- successors 1004 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3221_if_link/$entry
      -- 
    cp_elements(1003) <= cp_elements(1002);
    -- CP-element group 1004 transition  place  input  bypass 
    -- predecessors 1003 
    -- successors 2040 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3221_if_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3221_if_link/if_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi
      -- 
    if_choice_transition_12558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3221_branch_ack_1, ack => cp_elements(1004)); -- 
    -- CP-element group 1005 transition  bypass 
    -- predecessors 1002 
    -- successors 1006 
    -- members (1) 
      -- 	branch_block_stmt_1659/if_stmt_3221_else_link/$entry
      -- 
    cp_elements(1005) <= cp_elements(1002);
    -- CP-element group 1006 transition  place  input  bypass 
    -- predecessors 1005 
    -- successors 2083 
    -- members (3) 
      -- 	branch_block_stmt_1659/if_stmt_3221_else_link/$exit
      -- 	branch_block_stmt_1659/if_stmt_3221_else_link/else_choice_transition
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi
      -- 
    else_choice_transition_12562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3221_branch_ack_0, ack => cp_elements(1006)); -- 
    -- CP-element group 1007 fork  transition  bypass 
    -- predecessors 60 
    -- successors 1008 1009 1013 1014 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/$entry
      -- 
    cp_elements(1007) <= cp_elements(60);
    -- CP-element group 1008 transition  output  bypass 
    -- predecessors 1007 
    -- successors 1011 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Update/cr
      -- 
    cp_elements(1008) <= cp_elements(1007);
    cr_12584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1008), ack => ADD_u32_u32_3241_inst_req_1); -- 
    -- CP-element group 1009 transition  output  bypass 
    -- predecessors 1007 
    -- successors 1010 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_iNsTr_196_3238_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_iNsTr_196_3238_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_iNsTr_196_3238_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_iNsTr_196_3238_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Sample/rr
      -- 
    cp_elements(1009) <= cp_elements(1007);
    rr_12579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1009), ack => ADD_u32_u32_3241_inst_req_0); -- 
    -- CP-element group 1010 transition  input  bypass 
    -- predecessors 1009 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Sample/ra
      -- 
    ra_12580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3241_inst_ack_0, ack => cp_elements(1010)); -- 
    -- CP-element group 1011 transition  input  bypass 
    -- predecessors 1008 
    -- successors 1012 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/ADD_u32_u32_3241_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_tmp25x_xi_3244_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_tmp25x_xi_3244_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_tmp25x_xi_3244_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_tmp25x_xi_3244_update_completed_
      -- 
    ca_12585_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3241_inst_ack_1, ack => cp_elements(1011)); -- 
    -- CP-element group 1012 join  transition  output  bypass 
    -- predecessors 1011 1014 
    -- successors 1015 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Sample/rr
      -- 
    cp_element_group_1012: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1012"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1011) & cp_elements(1014);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1012), clk => clk, reset => reset); --
    end block;
    rr_12601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1012), ack => SUB_u32_u32_3246_inst_req_0); -- 
    -- CP-element group 1013 transition  output  bypass 
    -- predecessors 1007 
    -- successors 1016 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Update/cr
      -- 
    cp_elements(1013) <= cp_elements(1007);
    cr_12606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1013), ack => SUB_u32_u32_3246_inst_req_1); -- 
    -- CP-element group 1014 transition  bypass 
    -- predecessors 1007 
    -- successors 1012 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_xx_xlcssa_3245_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_xx_xlcssa_3245_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_xx_xlcssa_3245_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/R_xx_xlcssa_3245_update_completed_
      -- 
    cp_elements(1014) <= cp_elements(1007);
    -- CP-element group 1015 transition  input  bypass 
    -- predecessors 1012 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Sample/ra
      -- 
    ra_12602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3246_inst_ack_0, ack => cp_elements(1015)); -- 
    -- CP-element group 1016 transition  place  input  bypass 
    -- predecessors 1013 
    -- successors 2128 
    -- members (6) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3242_to_assign_stmt_3247/SUB_u32_u32_3246_Update/ca
      -- 
    ca_12607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_3246_inst_ack_1, ack => cp_elements(1016)); -- 
    -- CP-element group 1017 fork  transition  bypass 
    -- predecessors 61 
    -- successors 1018 1019 1022 1023 1026 1030 1031 1035 1038 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/$entry
      -- 
    cp_elements(1017) <= cp_elements(61);
    -- CP-element group 1018 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1021 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Update/cr
      -- 
    cp_elements(1018) <= cp_elements(1017);
    cr_12627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1018), ack => AND_u32_u32_3267_inst_req_1); -- 
    -- CP-element group 1019 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1020 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_tempx_x0x_xlcssax_xi_3264_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_tempx_x0x_xlcssax_xi_3264_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_tempx_x0x_xlcssax_xi_3264_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_tempx_x0x_xlcssax_xi_3264_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Sample/rr
      -- 
    cp_elements(1019) <= cp_elements(1017);
    rr_12622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1019), ack => AND_u32_u32_3267_inst_req_0); -- 
    -- CP-element group 1020 transition  input  bypass 
    -- predecessors 1019 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Sample/ra
      -- 
    ra_12623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3267_inst_ack_0, ack => cp_elements(1020)); -- 
    -- CP-element group 1021 transition  input  bypass 
    -- predecessors 1018 
    -- successors 1034 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/AND_u32_u32_3267_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_205_3288_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_205_3288_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_205_3288_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_205_3288_update_completed_
      -- 
    ca_12628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_3267_inst_ack_1, ack => cp_elements(1021)); -- 
    -- CP-element group 1022 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1025 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Update/cr
      -- 
    cp_elements(1022) <= cp_elements(1017);
    cr_12645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1022), ack => SHL_u32_u32_3273_inst_req_1); -- 
    -- CP-element group 1023 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1024 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_expx_x0x_xlcssax_xi_3270_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_expx_x0x_xlcssax_xi_3270_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_expx_x0x_xlcssax_xi_3270_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_expx_x0x_xlcssax_xi_3270_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Sample/rr
      -- 
    cp_elements(1023) <= cp_elements(1017);
    rr_12640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1023), ack => SHL_u32_u32_3273_inst_req_0); -- 
    -- CP-element group 1024 transition  input  bypass 
    -- predecessors 1023 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Sample/ra
      -- 
    ra_12641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3273_inst_ack_0, ack => cp_elements(1024)); -- 
    -- CP-element group 1025 transition  input  output  bypass 
    -- predecessors 1022 
    -- successors 1027 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/SHL_u32_u32_3273_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_206_3276_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_206_3276_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_206_3276_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_206_3276_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Sample/rr
      -- 
    ca_12646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_3273_inst_ack_1, ack => cp_elements(1025)); -- 
    rr_12658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1025), ack => ADD_u32_u32_3279_inst_req_0); -- 
    -- CP-element group 1026 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1028 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Update/cr
      -- 
    cp_elements(1026) <= cp_elements(1017);
    cr_12663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1026), ack => ADD_u32_u32_3279_inst_req_1); -- 
    -- CP-element group 1027 transition  input  bypass 
    -- predecessors 1025 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Sample/ra
      -- 
    ra_12659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3279_inst_ack_0, ack => cp_elements(1027)); -- 
    -- CP-element group 1028 transition  input  bypass 
    -- predecessors 1026 
    -- successors 1029 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/ADD_u32_u32_3279_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_207_3282_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_207_3282_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_207_3282_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_207_3282_update_completed_
      -- 
    ca_12664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_3279_inst_ack_1, ack => cp_elements(1028)); -- 
    -- CP-element group 1029 join  transition  output  bypass 
    -- predecessors 1028 1031 
    -- successors 1032 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Sample/rr
      -- 
    cp_element_group_1029: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1029"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1028) & cp_elements(1031);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1029), clk => clk, reset => reset); --
    end block;
    rr_12680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1029), ack => OR_u32_u32_3284_inst_req_0); -- 
    -- CP-element group 1030 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1033 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Update/cr
      -- 
    cp_elements(1030) <= cp_elements(1017);
    cr_12685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1030), ack => OR_u32_u32_3284_inst_req_1); -- 
    -- CP-element group 1031 transition  bypass 
    -- predecessors 1017 
    -- successors 1029 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_195_3283_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_195_3283_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_195_3283_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_195_3283_update_completed_
      -- 
    cp_elements(1031) <= cp_elements(1017);
    -- CP-element group 1032 transition  input  bypass 
    -- predecessors 1029 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Sample/ra
      -- 
    ra_12681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3284_inst_ack_0, ack => cp_elements(1032)); -- 
    -- CP-element group 1033 transition  input  bypass 
    -- predecessors 1030 
    -- successors 1034 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3284_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_208_3287_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_208_3287_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_208_3287_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_208_3287_update_completed_
      -- 
    ca_12686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3284_inst_ack_1, ack => cp_elements(1033)); -- 
    -- CP-element group 1034 join  transition  output  bypass 
    -- predecessors 1021 1033 
    -- successors 1036 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Sample/rr
      -- 
    cp_element_group_1034: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1034"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1021) & cp_elements(1033);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1034), clk => clk, reset => reset); --
    end block;
    rr_12702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1034), ack => OR_u32_u32_3289_inst_req_0); -- 
    -- CP-element group 1035 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1037 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Update/cr
      -- 
    cp_elements(1035) <= cp_elements(1017);
    cr_12707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1035), ack => OR_u32_u32_3289_inst_req_1); -- 
    -- CP-element group 1036 transition  input  bypass 
    -- predecessors 1034 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Sample/ra
      -- 
    ra_12703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3289_inst_ack_0, ack => cp_elements(1036)); -- 
    -- CP-element group 1037 transition  input  output  bypass 
    -- predecessors 1035 
    -- successors 1039 
    -- members (10) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_209_3292_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/OR_u32_u32_3289_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_209_3292_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_209_3292_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/R_iNsTr_209_3292_update_start_
      -- 
    ca_12708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_3289_inst_ack_1, ack => cp_elements(1037)); -- 
    rr_12720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1037), ack => type_cast_3293_inst_req_0); -- 
    -- CP-element group 1038 transition  output  bypass 
    -- predecessors 1017 
    -- successors 1040 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Update/cr
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_update_start_
      -- 
    cp_elements(1038) <= cp_elements(1017);
    cr_12725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1038), ack => type_cast_3293_inst_req_1); -- 
    -- CP-element group 1039 transition  input  bypass 
    -- predecessors 1037 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_sample_completed_
      -- 
    ra_12721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3293_inst_ack_0, ack => cp_elements(1039)); -- 
    -- CP-element group 1040 fork  transition  place  input  bypass 
    -- predecessors 1038 
    -- successors 2162 2164 
    -- members (11) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Update/ca
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3268_to_assign_stmt_3294/type_cast_3293_update_completed_
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/$entry
      -- 
    ca_12726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3293_inst_ack_1, ack => cp_elements(1040)); -- 
    -- CP-element group 1041 fork  transition  bypass 
    -- predecessors 2169 
    -- successors 1042 1043 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3307/$entry
      -- 
    cp_elements(1041) <= cp_elements(2169);
    -- CP-element group 1042 transition  output  bypass 
    -- predecessors 1041 
    -- successors 1044 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3307/R_iNsTr_173_3306_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3307/R_iNsTr_173_3306_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3307/R_iNsTr_173_3306_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3307/R_iNsTr_173_3306_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Sample/req
      -- 
    cp_elements(1042) <= cp_elements(1041);
    req_12741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1042), ack => WPIPE_out_data_3305_inst_req_0); -- 
    -- CP-element group 1043 transition  output  bypass 
    -- predecessors 1041 
    -- successors 1045 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Update/req
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Update/$entry
      -- 
    cp_elements(1043) <= cp_elements(1041);
    req_12746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1043), ack => WPIPE_out_data_3305_inst_req_1); -- 
    -- CP-element group 1044 transition  input  bypass 
    -- predecessors 1042 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Sample/ack
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Sample/$exit
      -- 
    ack_12742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3305_inst_ack_0, ack => cp_elements(1044)); -- 
    -- CP-element group 1045 transition  place  input  bypass 
    -- predecessors 1043 
    -- successors 1046 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3310__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3307__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3307/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Update/ack
      -- 	branch_block_stmt_1659/assign_stmt_3307/WPIPE_out_data_3305_Update/$exit
      -- 
    ack_12747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3305_inst_ack_1, ack => cp_elements(1045)); -- 
    -- CP-element group 1046 fork  transition  bypass 
    -- predecessors 1045 
    -- successors 1047 1048 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3310/$entry
      -- 
    cp_elements(1046) <= cp_elements(1045);
    -- CP-element group 1047 transition  output  bypass 
    -- predecessors 1046 
    -- successors 1049 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3310/R_iNsTr_67_3309_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3310/R_iNsTr_67_3309_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Sample/req
      -- 	branch_block_stmt_1659/assign_stmt_3310/R_iNsTr_67_3309_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3310/R_iNsTr_67_3309_sample_start_
      -- 
    cp_elements(1047) <= cp_elements(1046);
    req_12762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1047), ack => WPIPE_out_data_3308_inst_req_0); -- 
    -- CP-element group 1048 transition  output  bypass 
    -- predecessors 1046 
    -- successors 1050 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Update/req
      -- 
    cp_elements(1048) <= cp_elements(1046);
    req_12767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1048), ack => WPIPE_out_data_3308_inst_req_1); -- 
    -- CP-element group 1049 transition  input  bypass 
    -- predecessors 1047 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Sample/ack
      -- 
    ack_12763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3308_inst_ack_0, ack => cp_elements(1049)); -- 
    -- CP-element group 1050 transition  place  input  bypass 
    -- predecessors 1048 
    -- successors 1051 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3313__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3310__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3310/WPIPE_out_data_3308_Update/ack
      -- 	branch_block_stmt_1659/assign_stmt_3310/$exit
      -- 
    ack_12768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3308_inst_ack_1, ack => cp_elements(1050)); -- 
    -- CP-element group 1051 fork  transition  bypass 
    -- predecessors 1050 
    -- successors 1052 1053 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3313/$entry
      -- 
    cp_elements(1051) <= cp_elements(1050);
    -- CP-element group 1052 transition  output  bypass 
    -- predecessors 1051 
    -- successors 1054 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Sample/req
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3313/R_iNsTr_49_3312_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3313/R_iNsTr_49_3312_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3313/R_iNsTr_49_3312_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3313/R_iNsTr_49_3312_sample_completed_
      -- 
    cp_elements(1052) <= cp_elements(1051);
    req_12783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1052), ack => WPIPE_out_data_3311_inst_req_0); -- 
    -- CP-element group 1053 transition  output  bypass 
    -- predecessors 1051 
    -- successors 1055 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Update/req
      -- 
    cp_elements(1053) <= cp_elements(1051);
    req_12788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1053), ack => WPIPE_out_data_3311_inst_req_1); -- 
    -- CP-element group 1054 transition  input  bypass 
    -- predecessors 1052 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Sample/ack
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Sample/$exit
      -- 
    ack_12784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3311_inst_ack_0, ack => cp_elements(1054)); -- 
    -- CP-element group 1055 transition  place  input  bypass 
    -- predecessors 1053 
    -- successors 1056 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3313__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3316__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3313/WPIPE_out_data_3311_Update/ack
      -- 	branch_block_stmt_1659/assign_stmt_3313/$exit
      -- 
    ack_12789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3311_inst_ack_1, ack => cp_elements(1055)); -- 
    -- CP-element group 1056 fork  transition  bypass 
    -- predecessors 1055 
    -- successors 1057 1058 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3316/$entry
      -- 
    cp_elements(1056) <= cp_elements(1055);
    -- CP-element group 1057 transition  output  bypass 
    -- predecessors 1056 
    -- successors 1059 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3316/R_iNsTr_39_3315_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3316/R_iNsTr_39_3315_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3316/R_iNsTr_39_3315_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Sample/req
      -- 	branch_block_stmt_1659/assign_stmt_3316/R_iNsTr_39_3315_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Sample/$entry
      -- 
    cp_elements(1057) <= cp_elements(1056);
    req_12804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1057), ack => WPIPE_out_data_3314_inst_req_0); -- 
    -- CP-element group 1058 transition  output  bypass 
    -- predecessors 1056 
    -- successors 1060 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Update/req
      -- 
    cp_elements(1058) <= cp_elements(1056);
    req_12809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1058), ack => WPIPE_out_data_3314_inst_req_1); -- 
    -- CP-element group 1059 transition  input  bypass 
    -- predecessors 1057 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Sample/ack
      -- 
    ack_12805_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3314_inst_ack_0, ack => cp_elements(1059)); -- 
    -- CP-element group 1060 transition  place  input  bypass 
    -- predecessors 1058 
    -- successors 1061 
    -- members (6) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334__entry__
      -- 	branch_block_stmt_1659/assign_stmt_3316__exit__
      -- 	branch_block_stmt_1659/assign_stmt_3316/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Update/ack
      -- 	branch_block_stmt_1659/assign_stmt_3316/WPIPE_out_data_3314_Update/$exit
      -- 
    ack_12810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3314_inst_ack_1, ack => cp_elements(1060)); -- 
    -- CP-element group 1061 fork  transition  bypass 
    -- predecessors 1060 
    -- successors 1062 1063 1066 1067 1070 1071 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/$entry
      -- 
    cp_elements(1061) <= cp_elements(1060);
    -- CP-element group 1062 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1065 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Update/cr
      -- 
    cp_elements(1062) <= cp_elements(1061);
    cr_12830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1062), ack => MUL_f32_f32_3321_inst_req_1); -- 
    -- CP-element group 1063 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1064 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_20_3318_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Sample/rr
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_20_3318_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_20_3318_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_20_3318_sample_start_
      -- 
    cp_elements(1063) <= cp_elements(1061);
    rr_12825_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1063), ack => MUL_f32_f32_3321_inst_req_0); -- 
    -- CP-element group 1064 transition  input  bypass 
    -- predecessors 1063 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Sample/ra
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Sample/$exit
      -- 
    ra_12826_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3321_inst_ack_0, ack => cp_elements(1064)); -- 
    -- CP-element group 1065 transition  input  bypass 
    -- predecessors 1062 
    -- successors 1074 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3321_Update/ca
      -- 
    ca_12831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3321_inst_ack_1, ack => cp_elements(1065)); -- 
    -- CP-element group 1066 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1069 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Update/cr
      -- 
    cp_elements(1066) <= cp_elements(1061);
    cr_12848_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1066), ack => MUL_f32_f32_3327_inst_req_1); -- 
    -- CP-element group 1067 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1068 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_39_3324_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_39_3324_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_39_3324_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_39_3324_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Sample/rr
      -- 
    cp_elements(1067) <= cp_elements(1061);
    rr_12843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1067), ack => MUL_f32_f32_3327_inst_req_0); -- 
    -- CP-element group 1068 transition  input  bypass 
    -- predecessors 1067 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Sample/ra
      -- 
    ra_12844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3327_inst_ack_0, ack => cp_elements(1068)); -- 
    -- CP-element group 1069 transition  input  bypass 
    -- predecessors 1066 
    -- successors 1074 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3327_Update/ca
      -- 
    ca_12849_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3327_inst_ack_1, ack => cp_elements(1069)); -- 
    -- CP-element group 1070 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1073 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Update/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Update/cr
      -- 
    cp_elements(1070) <= cp_elements(1061);
    cr_12866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1070), ack => MUL_f32_f32_3333_inst_req_1); -- 
    -- CP-element group 1071 transition  output  bypass 
    -- predecessors 1061 
    -- successors 1072 
    -- members (7) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_69_3330_sample_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_69_3330_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_69_3330_update_start_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/R_iNsTr_69_3330_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Sample/$entry
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Sample/rr
      -- 
    cp_elements(1071) <= cp_elements(1061);
    rr_12861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1071), ack => MUL_f32_f32_3333_inst_req_0); -- 
    -- CP-element group 1072 transition  input  bypass 
    -- predecessors 1071 
    -- successors 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_sample_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Sample/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Sample/ra
      -- 
    ra_12862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3333_inst_ack_0, ack => cp_elements(1072)); -- 
    -- CP-element group 1073 transition  input  bypass 
    -- predecessors 1070 
    -- successors 1074 
    -- members (3) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_update_completed_
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Update/$exit
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/MUL_f32_f32_3333_Update/ca
      -- 
    ca_12867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_3333_inst_ack_1, ack => cp_elements(1073)); -- 
    -- CP-element group 1074 join  transition  bypass 
    -- predecessors 1065 1069 1073 
    -- successors 62 
    -- members (1) 
      -- 	branch_block_stmt_1659/assign_stmt_3322_to_assign_stmt_3334/$exit
      -- 
    cp_element_group_1074: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1074"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1065) & cp_elements(1069) & cp_elements(1073);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1074), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1075 fork  transition  bypass 
    -- predecessors 0 
    -- successors 1076 1080 1084 1088 1092 1096 1100 1104 
    -- members (1) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/$entry
      -- 
    cp_elements(1075) <= cp_elements(0);
    -- CP-element group 1076 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1077 1078 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/$entry
      -- 
    cp_elements(1076) <= cp_elements(1075);
    -- CP-element group 1077 transition  bypass 
    -- predecessors 1076 
    -- successors 1079 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/ra
      -- 
    cp_elements(1077) <= cp_elements(1076);
    -- CP-element group 1078 transition  bypass 
    -- predecessors 1076 
    -- successors 1079 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/ca
      -- 
    cp_elements(1078) <= cp_elements(1076);
    -- CP-element group 1079 join  transition  output  bypass 
    -- predecessors 1077 1078 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_req
      -- 
    cp_element_group_1079: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1079"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1077) & cp_elements(1078);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1079), clk => clk, reset => reset); --
    end block;
    phi_stmt_1697_req_12893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1079), ack => phi_stmt_1697_req_0); -- 
    -- CP-element group 1080 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1081 1082 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/$entry
      -- 
    cp_elements(1080) <= cp_elements(1075);
    -- CP-element group 1081 transition  bypass 
    -- predecessors 1080 
    -- successors 1083 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/ra
      -- 
    cp_elements(1081) <= cp_elements(1080);
    -- CP-element group 1082 transition  bypass 
    -- predecessors 1080 
    -- successors 1083 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/ca
      -- 
    cp_elements(1082) <= cp_elements(1080);
    -- CP-element group 1083 join  transition  output  bypass 
    -- predecessors 1081 1082 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_req
      -- 
    cp_element_group_1083: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1083"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1081) & cp_elements(1082);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1083), clk => clk, reset => reset); --
    end block;
    phi_stmt_1683_req_12916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1083), ack => phi_stmt_1683_req_0); -- 
    -- CP-element group 1084 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1085 1086 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/$entry
      -- 
    cp_elements(1084) <= cp_elements(1075);
    -- CP-element group 1085 transition  bypass 
    -- predecessors 1084 
    -- successors 1087 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/ra
      -- 
    cp_elements(1085) <= cp_elements(1084);
    -- CP-element group 1086 transition  bypass 
    -- predecessors 1084 
    -- successors 1087 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/ca
      -- 
    cp_elements(1086) <= cp_elements(1084);
    -- CP-element group 1087 join  transition  output  bypass 
    -- predecessors 1085 1086 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_req
      -- 
    cp_element_group_1087: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1087"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1085) & cp_elements(1086);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1087), clk => clk, reset => reset); --
    end block;
    phi_stmt_1704_req_12939_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1087), ack => phi_stmt_1704_req_0); -- 
    -- CP-element group 1088 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1089 1090 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/$entry
      -- 
    cp_elements(1088) <= cp_elements(1075);
    -- CP-element group 1089 transition  bypass 
    -- predecessors 1088 
    -- successors 1091 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/ra
      -- 
    cp_elements(1089) <= cp_elements(1088);
    -- CP-element group 1090 transition  bypass 
    -- predecessors 1088 
    -- successors 1091 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/ca
      -- 
    cp_elements(1090) <= cp_elements(1088);
    -- CP-element group 1091 join  transition  output  bypass 
    -- predecessors 1089 1090 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_req
      -- 
    cp_element_group_1091: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1091"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1089) & cp_elements(1090);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1091), clk => clk, reset => reset); --
    end block;
    phi_stmt_1676_req_12962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1091), ack => phi_stmt_1676_req_0); -- 
    -- CP-element group 1092 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1093 1094 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/$entry
      -- 
    cp_elements(1092) <= cp_elements(1075);
    -- CP-element group 1093 transition  bypass 
    -- predecessors 1092 
    -- successors 1095 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/ra
      -- 
    cp_elements(1093) <= cp_elements(1092);
    -- CP-element group 1094 transition  bypass 
    -- predecessors 1092 
    -- successors 1095 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/ca
      -- 
    cp_elements(1094) <= cp_elements(1092);
    -- CP-element group 1095 join  transition  output  bypass 
    -- predecessors 1093 1094 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_req
      -- 
    cp_element_group_1095: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1095"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1093) & cp_elements(1094);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1095), clk => clk, reset => reset); --
    end block;
    phi_stmt_1711_req_12985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1095), ack => phi_stmt_1711_req_0); -- 
    -- CP-element group 1096 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1097 1098 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/$entry
      -- 
    cp_elements(1096) <= cp_elements(1075);
    -- CP-element group 1097 transition  bypass 
    -- predecessors 1096 
    -- successors 1099 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/ra
      -- 
    cp_elements(1097) <= cp_elements(1096);
    -- CP-element group 1098 transition  bypass 
    -- predecessors 1096 
    -- successors 1099 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/ca
      -- 
    cp_elements(1098) <= cp_elements(1096);
    -- CP-element group 1099 join  transition  output  bypass 
    -- predecessors 1097 1098 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_req
      -- 
    cp_element_group_1099: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1099"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1097) & cp_elements(1098);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1099), clk => clk, reset => reset); --
    end block;
    phi_stmt_1669_req_13008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1099), ack => phi_stmt_1669_req_0); -- 
    -- CP-element group 1100 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1101 1102 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/$entry
      -- 
    cp_elements(1100) <= cp_elements(1075);
    -- CP-element group 1101 transition  bypass 
    -- predecessors 1100 
    -- successors 1103 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/ra
      -- 
    cp_elements(1101) <= cp_elements(1100);
    -- CP-element group 1102 transition  bypass 
    -- predecessors 1100 
    -- successors 1103 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/ca
      -- 
    cp_elements(1102) <= cp_elements(1100);
    -- CP-element group 1103 join  transition  output  bypass 
    -- predecessors 1101 1102 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_req
      -- 
    cp_element_group_1103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1101) & cp_elements(1102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1103), clk => clk, reset => reset); --
    end block;
    phi_stmt_1690_req_13031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1103), ack => phi_stmt_1690_req_0); -- 
    -- CP-element group 1104 fork  transition  bypass 
    -- predecessors 1075 
    -- successors 1105 1106 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/$entry
      -- 
    cp_elements(1104) <= cp_elements(1075);
    -- CP-element group 1105 transition  bypass 
    -- predecessors 1104 
    -- successors 1107 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/ra
      -- 
    cp_elements(1105) <= cp_elements(1104);
    -- CP-element group 1106 transition  bypass 
    -- predecessors 1104 
    -- successors 1107 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/ca
      -- 
    cp_elements(1106) <= cp_elements(1104);
    -- CP-element group 1107 join  transition  output  bypass 
    -- predecessors 1105 1106 
    -- successors 1108 
    -- members (5) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_req
      -- 
    cp_element_group_1107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1105) & cp_elements(1106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1107), clk => clk, reset => reset); --
    end block;
    phi_stmt_1662_req_13054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1107), ack => phi_stmt_1662_req_0); -- 
    -- CP-element group 1108 join  transition  bypass 
    -- predecessors 1079 1083 1087 1091 1095 1099 1103 1107 
    -- successors 1159 
    -- members (1) 
      -- 	branch_block_stmt_1659/bb_0_bb_1_PhiReq/$exit
      -- 
    cp_element_group_1108: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1108"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= cp_elements(1079) & cp_elements(1083) & cp_elements(1087) & cp_elements(1091) & cp_elements(1095) & cp_elements(1099) & cp_elements(1103) & cp_elements(1107);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1109 fork  transition  bypass 
    -- predecessors 62 
    -- successors 1110 1116 1122 1128 1134 1140 1146 1152 
    -- members (1) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/$entry
      -- 
    cp_elements(1109) <= cp_elements(62);
    -- CP-element group 1110 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1111 1113 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/$entry
      -- 
    cp_elements(1110) <= cp_elements(1109);
    -- CP-element group 1111 transition  output  bypass 
    -- predecessors 1110 
    -- successors 1112 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/rr
      -- 
    cp_elements(1111) <= cp_elements(1110);
    rr_13073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1111), ack => type_cast_1703_inst_req_0); -- 
    -- CP-element group 1112 transition  input  bypass 
    -- predecessors 1111 
    -- successors 1115 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Sample/ra
      -- 
    ra_13074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1703_inst_ack_0, ack => cp_elements(1112)); -- 
    -- CP-element group 1113 transition  output  bypass 
    -- predecessors 1110 
    -- successors 1114 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/cr
      -- 
    cp_elements(1113) <= cp_elements(1110);
    cr_13078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1113), ack => type_cast_1703_inst_req_1); -- 
    -- CP-element group 1114 transition  input  bypass 
    -- predecessors 1113 
    -- successors 1115 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/Update/ca
      -- 
    ca_13079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1703_inst_ack_1, ack => cp_elements(1114)); -- 
    -- CP-element group 1115 join  transition  output  bypass 
    -- predecessors 1112 1114 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_sources/type_cast_1703/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1697/phi_stmt_1697_req
      -- 
    cp_element_group_1115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1112) & cp_elements(1114);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1115), clk => clk, reset => reset); --
    end block;
    phi_stmt_1697_req_13080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1115), ack => phi_stmt_1697_req_1); -- 
    -- CP-element group 1116 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1117 1119 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/$entry
      -- 
    cp_elements(1116) <= cp_elements(1109);
    -- CP-element group 1117 transition  output  bypass 
    -- predecessors 1116 
    -- successors 1118 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/rr
      -- 
    cp_elements(1117) <= cp_elements(1116);
    rr_13096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1117), ack => type_cast_1689_inst_req_0); -- 
    -- CP-element group 1118 transition  input  bypass 
    -- predecessors 1117 
    -- successors 1121 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Sample/ra
      -- 
    ra_13097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_0, ack => cp_elements(1118)); -- 
    -- CP-element group 1119 transition  output  bypass 
    -- predecessors 1116 
    -- successors 1120 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/cr
      -- 
    cp_elements(1119) <= cp_elements(1116);
    cr_13101_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1119), ack => type_cast_1689_inst_req_1); -- 
    -- CP-element group 1120 transition  input  bypass 
    -- predecessors 1119 
    -- successors 1121 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/Update/ca
      -- 
    ca_13102_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_1, ack => cp_elements(1120)); -- 
    -- CP-element group 1121 join  transition  output  bypass 
    -- predecessors 1118 1120 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_sources/type_cast_1689/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1683/phi_stmt_1683_req
      -- 
    cp_element_group_1121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1118) & cp_elements(1120);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1121), clk => clk, reset => reset); --
    end block;
    phi_stmt_1683_req_13103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1121), ack => phi_stmt_1683_req_1); -- 
    -- CP-element group 1122 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1123 1125 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/$entry
      -- 
    cp_elements(1122) <= cp_elements(1109);
    -- CP-element group 1123 transition  output  bypass 
    -- predecessors 1122 
    -- successors 1124 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/rr
      -- 
    cp_elements(1123) <= cp_elements(1122);
    rr_13119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1123), ack => type_cast_1710_inst_req_0); -- 
    -- CP-element group 1124 transition  input  bypass 
    -- predecessors 1123 
    -- successors 1127 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Sample/ra
      -- 
    ra_13120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_0, ack => cp_elements(1124)); -- 
    -- CP-element group 1125 transition  output  bypass 
    -- predecessors 1122 
    -- successors 1126 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/cr
      -- 
    cp_elements(1125) <= cp_elements(1122);
    cr_13124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1125), ack => type_cast_1710_inst_req_1); -- 
    -- CP-element group 1126 transition  input  bypass 
    -- predecessors 1125 
    -- successors 1127 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/Update/ca
      -- 
    ca_13125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_1, ack => cp_elements(1126)); -- 
    -- CP-element group 1127 join  transition  output  bypass 
    -- predecessors 1124 1126 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_sources/type_cast_1710/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1704/phi_stmt_1704_req
      -- 
    cp_element_group_1127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1124) & cp_elements(1126);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1127), clk => clk, reset => reset); --
    end block;
    phi_stmt_1704_req_13126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1127), ack => phi_stmt_1704_req_1); -- 
    -- CP-element group 1128 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1129 1131 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/$entry
      -- 
    cp_elements(1128) <= cp_elements(1109);
    -- CP-element group 1129 transition  output  bypass 
    -- predecessors 1128 
    -- successors 1130 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/rr
      -- 
    cp_elements(1129) <= cp_elements(1128);
    rr_13142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1129), ack => type_cast_1682_inst_req_0); -- 
    -- CP-element group 1130 transition  input  bypass 
    -- predecessors 1129 
    -- successors 1133 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Sample/ra
      -- 
    ra_13143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1682_inst_ack_0, ack => cp_elements(1130)); -- 
    -- CP-element group 1131 transition  output  bypass 
    -- predecessors 1128 
    -- successors 1132 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/cr
      -- 
    cp_elements(1131) <= cp_elements(1128);
    cr_13147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1131), ack => type_cast_1682_inst_req_1); -- 
    -- CP-element group 1132 transition  input  bypass 
    -- predecessors 1131 
    -- successors 1133 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/Update/ca
      -- 
    ca_13148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1682_inst_ack_1, ack => cp_elements(1132)); -- 
    -- CP-element group 1133 join  transition  output  bypass 
    -- predecessors 1130 1132 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_sources/type_cast_1682/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1676/phi_stmt_1676_req
      -- 
    cp_element_group_1133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1130) & cp_elements(1132);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1133), clk => clk, reset => reset); --
    end block;
    phi_stmt_1676_req_13149_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1133), ack => phi_stmt_1676_req_1); -- 
    -- CP-element group 1134 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1135 1137 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/$entry
      -- 
    cp_elements(1134) <= cp_elements(1109);
    -- CP-element group 1135 transition  output  bypass 
    -- predecessors 1134 
    -- successors 1136 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/rr
      -- 
    cp_elements(1135) <= cp_elements(1134);
    rr_13165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1135), ack => type_cast_1717_inst_req_0); -- 
    -- CP-element group 1136 transition  input  bypass 
    -- predecessors 1135 
    -- successors 1139 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Sample/ra
      -- 
    ra_13166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_0, ack => cp_elements(1136)); -- 
    -- CP-element group 1137 transition  output  bypass 
    -- predecessors 1134 
    -- successors 1138 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/cr
      -- 
    cp_elements(1137) <= cp_elements(1134);
    cr_13170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1137), ack => type_cast_1717_inst_req_1); -- 
    -- CP-element group 1138 transition  input  bypass 
    -- predecessors 1137 
    -- successors 1139 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/Update/ca
      -- 
    ca_13171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_1, ack => cp_elements(1138)); -- 
    -- CP-element group 1139 join  transition  output  bypass 
    -- predecessors 1136 1138 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_sources/type_cast_1717/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1711/phi_stmt_1711_req
      -- 
    cp_element_group_1139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1136) & cp_elements(1138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1139), clk => clk, reset => reset); --
    end block;
    phi_stmt_1711_req_13172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1139), ack => phi_stmt_1711_req_1); -- 
    -- CP-element group 1140 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1141 1143 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/$entry
      -- 
    cp_elements(1140) <= cp_elements(1109);
    -- CP-element group 1141 transition  output  bypass 
    -- predecessors 1140 
    -- successors 1142 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/rr
      -- 
    cp_elements(1141) <= cp_elements(1140);
    rr_13188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1141), ack => type_cast_1675_inst_req_0); -- 
    -- CP-element group 1142 transition  input  bypass 
    -- predecessors 1141 
    -- successors 1145 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Sample/ra
      -- 
    ra_13189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_0, ack => cp_elements(1142)); -- 
    -- CP-element group 1143 transition  output  bypass 
    -- predecessors 1140 
    -- successors 1144 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/cr
      -- 
    cp_elements(1143) <= cp_elements(1140);
    cr_13193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1143), ack => type_cast_1675_inst_req_1); -- 
    -- CP-element group 1144 transition  input  bypass 
    -- predecessors 1143 
    -- successors 1145 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/Update/ca
      -- 
    ca_13194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_1, ack => cp_elements(1144)); -- 
    -- CP-element group 1145 join  transition  output  bypass 
    -- predecessors 1142 1144 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1675/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1669/phi_stmt_1669_req
      -- 
    cp_element_group_1145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1142) & cp_elements(1144);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1145), clk => clk, reset => reset); --
    end block;
    phi_stmt_1669_req_13195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1145), ack => phi_stmt_1669_req_1); -- 
    -- CP-element group 1146 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1147 1149 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/$entry
      -- 
    cp_elements(1146) <= cp_elements(1109);
    -- CP-element group 1147 transition  output  bypass 
    -- predecessors 1146 
    -- successors 1148 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/rr
      -- 
    cp_elements(1147) <= cp_elements(1146);
    rr_13211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1147), ack => type_cast_1696_inst_req_0); -- 
    -- CP-element group 1148 transition  input  bypass 
    -- predecessors 1147 
    -- successors 1151 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Sample/ra
      -- 
    ra_13212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1696_inst_ack_0, ack => cp_elements(1148)); -- 
    -- CP-element group 1149 transition  output  bypass 
    -- predecessors 1146 
    -- successors 1150 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/cr
      -- 
    cp_elements(1149) <= cp_elements(1146);
    cr_13216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1149), ack => type_cast_1696_inst_req_1); -- 
    -- CP-element group 1150 transition  input  bypass 
    -- predecessors 1149 
    -- successors 1151 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/Update/ca
      -- 
    ca_13217_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1696_inst_ack_1, ack => cp_elements(1150)); -- 
    -- CP-element group 1151 join  transition  output  bypass 
    -- predecessors 1148 1150 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1690/phi_stmt_1690_req
      -- 
    cp_element_group_1151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1148) & cp_elements(1150);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1151), clk => clk, reset => reset); --
    end block;
    phi_stmt_1690_req_13218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1151), ack => phi_stmt_1690_req_1); -- 
    -- CP-element group 1152 fork  transition  bypass 
    -- predecessors 1109 
    -- successors 1153 1155 
    -- members (4) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/$entry
      -- 
    cp_elements(1152) <= cp_elements(1109);
    -- CP-element group 1153 transition  output  bypass 
    -- predecessors 1152 
    -- successors 1154 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/rr
      -- 
    cp_elements(1153) <= cp_elements(1152);
    rr_13234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1153), ack => type_cast_1668_inst_req_0); -- 
    -- CP-element group 1154 transition  input  bypass 
    -- predecessors 1153 
    -- successors 1157 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Sample/ra
      -- 
    ra_13235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_0, ack => cp_elements(1154)); -- 
    -- CP-element group 1155 transition  output  bypass 
    -- predecessors 1152 
    -- successors 1156 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/cr
      -- 
    cp_elements(1155) <= cp_elements(1152);
    cr_13239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1155), ack => type_cast_1668_inst_req_1); -- 
    -- CP-element group 1156 transition  input  bypass 
    -- predecessors 1155 
    -- successors 1157 
    -- members (2) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/Update/ca
      -- 
    ca_13240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_1, ack => cp_elements(1156)); -- 
    -- CP-element group 1157 join  transition  output  bypass 
    -- predecessors 1154 1156 
    -- successors 1158 
    -- members (5) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1668/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/phi_stmt_1662/phi_stmt_1662_req
      -- 
    cp_element_group_1157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1154) & cp_elements(1156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1157), clk => clk, reset => reset); --
    end block;
    phi_stmt_1662_req_13241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1157), ack => phi_stmt_1662_req_1); -- 
    -- CP-element group 1158 join  transition  bypass 
    -- predecessors 1115 1121 1127 1133 1139 1145 1151 1157 
    -- successors 1159 
    -- members (1) 
      -- 	branch_block_stmt_1659/fdiv32x_xexit_bb_1_PhiReq/$exit
      -- 
    cp_element_group_1158: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1158"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= cp_elements(1115) & cp_elements(1121) & cp_elements(1127) & cp_elements(1133) & cp_elements(1139) & cp_elements(1145) & cp_elements(1151) & cp_elements(1157);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1159 merge  place  bypass 
    -- predecessors 1108 1158 
    -- successors 1160 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiReqMerge
      -- 
    cp_elements(1159) <= OrReduce(cp_elements(1108) & cp_elements(1158));
    -- CP-element group 1160 fork  transition  bypass 
    -- predecessors 1159 
    -- successors 1161 1162 1163 1164 1165 1166 1167 1168 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/$entry
      -- 
    cp_elements(1160) <= cp_elements(1159);
    -- CP-element group 1161 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1662_ack
      -- 
    phi_stmt_1662_ack_13246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1662_ack_0, ack => cp_elements(1161)); -- 
    -- CP-element group 1162 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1669_ack
      -- 
    phi_stmt_1669_ack_13247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1669_ack_0, ack => cp_elements(1162)); -- 
    -- CP-element group 1163 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1676_ack
      -- 
    phi_stmt_1676_ack_13248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1676_ack_0, ack => cp_elements(1163)); -- 
    -- CP-element group 1164 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1683_ack
      -- 
    phi_stmt_1683_ack_13249_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1683_ack_0, ack => cp_elements(1164)); -- 
    -- CP-element group 1165 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1690_ack
      -- 
    phi_stmt_1690_ack_13250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1690_ack_0, ack => cp_elements(1165)); -- 
    -- CP-element group 1166 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1697_ack
      -- 
    phi_stmt_1697_ack_13251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1697_ack_0, ack => cp_elements(1166)); -- 
    -- CP-element group 1167 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1704_ack
      -- 
    phi_stmt_1704_ack_13252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1704_ack_0, ack => cp_elements(1167)); -- 
    -- CP-element group 1168 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/phi_stmt_1711_ack
      -- 
    phi_stmt_1711_ack_13253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1711_ack_0, ack => cp_elements(1168)); -- 
    -- CP-element group 1169 join  transition  bypass 
    -- predecessors 1161 1162 1163 1164 1165 1166 1167 1168 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1661_PhiAck/$exit
      -- 
    cp_element_group_1169: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1169"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= cp_elements(1161) & cp_elements(1162) & cp_elements(1163) & cp_elements(1164) & cp_elements(1165) & cp_elements(1166) & cp_elements(1167) & cp_elements(1168);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1170 fork  transition  bypass 
    -- predecessors 112 
    -- successors 1171 1173 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$entry
      -- 
    cp_elements(1170) <= cp_elements(112);
    -- CP-element group 1171 transition  output  bypass 
    -- predecessors 1170 
    -- successors 1172 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/rr
      -- 
    cp_elements(1171) <= cp_elements(1170);
    rr_13304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1171), ack => type_cast_1794_inst_req_0); -- 
    -- CP-element group 1172 transition  input  bypass 
    -- predecessors 1171 
    -- successors 1175 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/ra
      -- 
    ra_13305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1794_inst_ack_0, ack => cp_elements(1172)); -- 
    -- CP-element group 1173 transition  output  bypass 
    -- predecessors 1170 
    -- successors 1174 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/cr
      -- 
    cp_elements(1173) <= cp_elements(1170);
    cr_13309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1173), ack => type_cast_1794_inst_req_1); -- 
    -- CP-element group 1174 transition  input  bypass 
    -- predecessors 1173 
    -- successors 1175 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/ca
      -- 
    ca_13310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1794_inst_ack_1, ack => cp_elements(1174)); -- 
    -- CP-element group 1175 join  transition  bypass 
    -- predecessors 1172 1174 
    -- successors 1184 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$exit
      -- 
    cp_element_group_1175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1172) & cp_elements(1174);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1176 fork  transition  bypass 
    -- predecessors 112 
    -- successors 1177 1178 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$entry
      -- 
    cp_elements(1176) <= cp_elements(112);
    -- CP-element group 1177 transition  bypass 
    -- predecessors 1176 
    -- successors 1179 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/ra
      -- 
    cp_elements(1177) <= cp_elements(1176);
    -- CP-element group 1178 transition  bypass 
    -- predecessors 1176 
    -- successors 1179 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/ca
      -- 
    cp_elements(1178) <= cp_elements(1176);
    -- CP-element group 1179 join  transition  bypass 
    -- predecessors 1177 1178 
    -- successors 1184 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$exit
      -- 
    cp_element_group_1179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1177) & cp_elements(1178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1180 fork  transition  bypass 
    -- predecessors 112 
    -- successors 1181 1182 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$entry
      -- 
    cp_elements(1180) <= cp_elements(112);
    -- CP-element group 1181 transition  bypass 
    -- predecessors 1180 
    -- successors 1183 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/ra
      -- 
    cp_elements(1181) <= cp_elements(1180);
    -- CP-element group 1182 transition  bypass 
    -- predecessors 1180 
    -- successors 1183 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/ca
      -- 
    cp_elements(1182) <= cp_elements(1180);
    -- CP-element group 1183 join  transition  bypass 
    -- predecessors 1181 1182 
    -- successors 1184 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$exit
      -- 
    cp_element_group_1183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1181) & cp_elements(1182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1184 join  transition  output  bypass 
    -- predecessors 1175 1179 1183 
    -- successors 1215 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$exit
      -- 	branch_block_stmt_1659/bb_2_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_req
      -- 
    cp_element_group_1184: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1184"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1175) & cp_elements(1179) & cp_elements(1183);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1184), clk => clk, reset => reset); --
    end block;
    phi_stmt_1791_req_13343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1184), ack => phi_stmt_1791_req_0); -- 
    -- CP-element group 1185 fork  transition  bypass 
    -- predecessors 126 
    -- successors 1186 1187 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$entry
      -- 
    cp_elements(1185) <= cp_elements(126);
    -- CP-element group 1186 transition  bypass 
    -- predecessors 1185 
    -- successors 1188 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/ra
      -- 
    cp_elements(1186) <= cp_elements(1185);
    -- CP-element group 1187 transition  bypass 
    -- predecessors 1185 
    -- successors 1188 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/ca
      -- 
    cp_elements(1187) <= cp_elements(1185);
    -- CP-element group 1188 join  transition  bypass 
    -- predecessors 1186 1187 
    -- successors 1199 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$exit
      -- 
    cp_element_group_1188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1186) & cp_elements(1187);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1189 fork  transition  bypass 
    -- predecessors 126 
    -- successors 1190 1191 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$entry
      -- 
    cp_elements(1189) <= cp_elements(126);
    -- CP-element group 1190 transition  bypass 
    -- predecessors 1189 
    -- successors 1192 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/ra
      -- 
    cp_elements(1190) <= cp_elements(1189);
    -- CP-element group 1191 transition  bypass 
    -- predecessors 1189 
    -- successors 1192 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/ca
      -- 
    cp_elements(1191) <= cp_elements(1189);
    -- CP-element group 1192 join  transition  bypass 
    -- predecessors 1190 1191 
    -- successors 1199 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$exit
      -- 
    cp_element_group_1192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1190) & cp_elements(1191);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1193 fork  transition  bypass 
    -- predecessors 126 
    -- successors 1194 1196 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$entry
      -- 
    cp_elements(1193) <= cp_elements(126);
    -- CP-element group 1194 transition  output  bypass 
    -- predecessors 1193 
    -- successors 1195 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/rr
      -- 
    cp_elements(1194) <= cp_elements(1193);
    rr_13394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1194), ack => type_cast_1798_inst_req_0); -- 
    -- CP-element group 1195 transition  input  bypass 
    -- predecessors 1194 
    -- successors 1198 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/ra
      -- 
    ra_13395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1798_inst_ack_0, ack => cp_elements(1195)); -- 
    -- CP-element group 1196 transition  output  bypass 
    -- predecessors 1193 
    -- successors 1197 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/cr
      -- 
    cp_elements(1196) <= cp_elements(1193);
    cr_13399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1196), ack => type_cast_1798_inst_req_1); -- 
    -- CP-element group 1197 transition  input  bypass 
    -- predecessors 1196 
    -- successors 1198 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/ca
      -- 
    ca_13400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1798_inst_ack_1, ack => cp_elements(1197)); -- 
    -- CP-element group 1198 join  transition  bypass 
    -- predecessors 1195 1197 
    -- successors 1199 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$exit
      -- 
    cp_element_group_1198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1195) & cp_elements(1197);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1199 join  transition  output  bypass 
    -- predecessors 1188 1192 1198 
    -- successors 1215 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$exit
      -- 	branch_block_stmt_1659/bb_3_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_req
      -- 
    cp_element_group_1199: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1199"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1188) & cp_elements(1192) & cp_elements(1198);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1199), clk => clk, reset => reset); --
    end block;
    phi_stmt_1791_req_13401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1199), ack => phi_stmt_1791_req_2); -- 
    -- CP-element group 1200 fork  transition  bypass 
    -- predecessors 137 
    -- successors 1201 1202 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$entry
      -- 
    cp_elements(1200) <= cp_elements(137);
    -- CP-element group 1201 transition  bypass 
    -- predecessors 1200 
    -- successors 1203 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Sample/ra
      -- 
    cp_elements(1201) <= cp_elements(1200);
    -- CP-element group 1202 transition  bypass 
    -- predecessors 1200 
    -- successors 1203 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/Update/ca
      -- 
    cp_elements(1202) <= cp_elements(1200);
    -- CP-element group 1203 join  transition  bypass 
    -- predecessors 1201 1202 
    -- successors 1214 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1794/SplitProtocol/$exit
      -- 
    cp_element_group_1203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1201) & cp_elements(1202);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1204 fork  transition  bypass 
    -- predecessors 137 
    -- successors 1205 1207 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$entry
      -- 
    cp_elements(1204) <= cp_elements(137);
    -- CP-element group 1205 transition  output  bypass 
    -- predecessors 1204 
    -- successors 1206 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/rr
      -- 
    cp_elements(1205) <= cp_elements(1204);
    rr_13436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1205), ack => type_cast_1796_inst_req_0); -- 
    -- CP-element group 1206 transition  input  bypass 
    -- predecessors 1205 
    -- successors 1209 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Sample/ra
      -- 
    ra_13437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_0, ack => cp_elements(1206)); -- 
    -- CP-element group 1207 transition  output  bypass 
    -- predecessors 1204 
    -- successors 1208 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/cr
      -- 
    cp_elements(1207) <= cp_elements(1204);
    cr_13441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1207), ack => type_cast_1796_inst_req_1); -- 
    -- CP-element group 1208 transition  input  bypass 
    -- predecessors 1207 
    -- successors 1209 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/Update/ca
      -- 
    ca_13442_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_1, ack => cp_elements(1208)); -- 
    -- CP-element group 1209 join  transition  bypass 
    -- predecessors 1206 1208 
    -- successors 1214 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1796/SplitProtocol/$exit
      -- 
    cp_element_group_1209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1206) & cp_elements(1208);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1210 fork  transition  bypass 
    -- predecessors 137 
    -- successors 1211 1212 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$entry
      -- 
    cp_elements(1210) <= cp_elements(137);
    -- CP-element group 1211 transition  bypass 
    -- predecessors 1210 
    -- successors 1213 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Sample/ra
      -- 
    cp_elements(1211) <= cp_elements(1210);
    -- CP-element group 1212 transition  bypass 
    -- predecessors 1210 
    -- successors 1213 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/Update/ca
      -- 
    cp_elements(1212) <= cp_elements(1210);
    -- CP-element group 1213 join  transition  bypass 
    -- predecessors 1211 1212 
    -- successors 1214 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/type_cast_1798/SplitProtocol/$exit
      -- 
    cp_element_group_1213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1211) & cp_elements(1212);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1214 join  transition  output  bypass 
    -- predecessors 1203 1209 1213 
    -- successors 1215 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_sources/$exit
      -- 	branch_block_stmt_1659/bb_4_bb_5_PhiReq/phi_stmt_1791/phi_stmt_1791_req
      -- 
    cp_element_group_1214: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1214"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= cp_elements(1203) & cp_elements(1209) & cp_elements(1213);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1214), clk => clk, reset => reset); --
    end block;
    phi_stmt_1791_req_13459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1214), ack => phi_stmt_1791_req_1); -- 
    -- CP-element group 1215 merge  place  bypass 
    -- predecessors 1184 1199 1214 
    -- successors 1216 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1790_PhiReqMerge
      -- 
    cp_elements(1215) <= OrReduce(cp_elements(1184) & cp_elements(1199) & cp_elements(1214));
    -- CP-element group 1216 transition  bypass 
    -- predecessors 1215 
    -- successors 1217 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1790_PhiAck/$entry
      -- 
    cp_elements(1216) <= cp_elements(1215);
    -- CP-element group 1217 transition  place  input  bypass 
    -- predecessors 1216 
    -- successors 138 
    -- members (4) 
      -- 	branch_block_stmt_1659/merge_stmt_1790__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1805_to_assign_stmt_1841__entry__
      -- 	branch_block_stmt_1659/merge_stmt_1790_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1790_PhiAck/phi_stmt_1791_ack
      -- 
    phi_stmt_1791_ack_13464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1791_ack_0, ack => cp_elements(1217)); -- 
    -- CP-element group 1218 transition  bypass 
    -- predecessors 176 
    -- successors 1220 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/ra
      -- 
    cp_elements(1218) <= cp_elements(176);
    -- CP-element group 1219 transition  bypass 
    -- predecessors 176 
    -- successors 1220 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/ca
      -- 
    cp_elements(1219) <= cp_elements(176);
    -- CP-element group 1220 join  transition  output  bypass 
    -- predecessors 1218 1219 
    -- successors 1229 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_5_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_req
      -- 
    cp_element_group_1220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1218) & cp_elements(1219);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1220), clk => clk, reset => reset); --
    end block;
    phi_stmt_1864_req_13514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1220), ack => phi_stmt_1864_req_1); -- 
    -- CP-element group 1221 transition  bypass 
    -- predecessors 188 
    -- successors 1223 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/ra
      -- 
    cp_elements(1221) <= cp_elements(188);
    -- CP-element group 1222 transition  bypass 
    -- predecessors 188 
    -- successors 1223 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/ca
      -- 
    cp_elements(1222) <= cp_elements(188);
    -- CP-element group 1223 join  transition  output  bypass 
    -- predecessors 1221 1222 
    -- successors 1229 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_6_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_req
      -- 
    cp_element_group_1223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1221) & cp_elements(1222);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1223), clk => clk, reset => reset); --
    end block;
    phi_stmt_1864_req_13540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1223), ack => phi_stmt_1864_req_2); -- 
    -- CP-element group 1224 transition  output  bypass 
    -- predecessors 6 
    -- successors 1225 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/rr
      -- 
    cp_elements(1224) <= cp_elements(6);
    rr_13559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1224), ack => type_cast_1867_inst_req_0); -- 
    -- CP-element group 1225 transition  input  bypass 
    -- predecessors 1224 
    -- successors 1228 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Sample/ra
      -- 
    ra_13560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_0, ack => cp_elements(1225)); -- 
    -- CP-element group 1226 transition  output  bypass 
    -- predecessors 6 
    -- successors 1227 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/cr
      -- 
    cp_elements(1226) <= cp_elements(6);
    cr_13564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1226), ack => type_cast_1867_inst_req_1); -- 
    -- CP-element group 1227 transition  input  bypass 
    -- predecessors 1226 
    -- successors 1228 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/Update/ca
      -- 
    ca_13565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_1, ack => cp_elements(1227)); -- 
    -- CP-element group 1228 join  transition  output  bypass 
    -- predecessors 1225 1227 
    -- successors 1229 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_sources/type_cast_1867/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_7_bb_8_PhiReq/phi_stmt_1864/phi_stmt_1864_req
      -- 
    cp_element_group_1228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1225) & cp_elements(1227);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1228), clk => clk, reset => reset); --
    end block;
    phi_stmt_1864_req_13566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1228), ack => phi_stmt_1864_req_0); -- 
    -- CP-element group 1229 merge  place  bypass 
    -- predecessors 1220 1223 1228 
    -- successors 1230 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1863_PhiReqMerge
      -- 
    cp_elements(1229) <= OrReduce(cp_elements(1220) & cp_elements(1223) & cp_elements(1228));
    -- CP-element group 1230 transition  bypass 
    -- predecessors 1229 
    -- successors 1231 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1863_PhiAck/$entry
      -- 
    cp_elements(1230) <= cp_elements(1229);
    -- CP-element group 1231 transition  place  input  bypass 
    -- predecessors 1230 
    -- successors 191 
    -- members (4) 
      -- 	branch_block_stmt_1659/merge_stmt_1863__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1880_to_assign_stmt_1891__entry__
      -- 	branch_block_stmt_1659/merge_stmt_1863_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1863_PhiAck/phi_stmt_1864_ack
      -- 
    phi_stmt_1864_ack_13571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1864_ack_0, ack => cp_elements(1231)); -- 
    -- CP-element group 1232 transition  output  bypass 
    -- predecessors 227 
    -- successors 1233 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/rr
      -- 
    cp_elements(1232) <= cp_elements(227);
    rr_13614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1232), ack => type_cast_1923_inst_req_0); -- 
    -- CP-element group 1233 transition  input  bypass 
    -- predecessors 1232 
    -- successors 1236 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/ra
      -- 
    ra_13615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_0, ack => cp_elements(1233)); -- 
    -- CP-element group 1234 transition  output  bypass 
    -- predecessors 227 
    -- successors 1235 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/cr
      -- 
    cp_elements(1234) <= cp_elements(227);
    cr_13619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1234), ack => type_cast_1923_inst_req_1); -- 
    -- CP-element group 1235 transition  input  bypass 
    -- predecessors 1234 
    -- successors 1236 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/ca
      -- 
    ca_13620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_1, ack => cp_elements(1235)); -- 
    -- CP-element group 1236 join  transition  output  bypass 
    -- predecessors 1233 1235 
    -- successors 1243 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_10_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_req
      -- 
    cp_element_group_1236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1233) & cp_elements(1235);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1236), clk => clk, reset => reset); --
    end block;
    phi_stmt_1920_req_13621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1236), ack => phi_stmt_1920_req_0); -- 
    -- CP-element group 1237 transition  bypass 
    -- predecessors 208 
    -- successors 1239 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/ra
      -- 
    cp_elements(1237) <= cp_elements(208);
    -- CP-element group 1238 transition  bypass 
    -- predecessors 208 
    -- successors 1239 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/ca
      -- 
    cp_elements(1238) <= cp_elements(208);
    -- CP-element group 1239 join  transition  output  bypass 
    -- predecessors 1237 1238 
    -- successors 1243 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_8_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_req
      -- 
    cp_element_group_1239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1237) & cp_elements(1238);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1239), clk => clk, reset => reset); --
    end block;
    phi_stmt_1920_req_13647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1239), ack => phi_stmt_1920_req_1); -- 
    -- CP-element group 1240 transition  bypass 
    -- predecessors 220 
    -- successors 1242 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Sample/ra
      -- 
    cp_elements(1240) <= cp_elements(220);
    -- CP-element group 1241 transition  bypass 
    -- predecessors 220 
    -- successors 1242 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/Update/ca
      -- 
    cp_elements(1241) <= cp_elements(220);
    -- CP-element group 1242 join  transition  output  bypass 
    -- predecessors 1240 1241 
    -- successors 1243 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_sources/type_cast_1923/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_9_bb_11_PhiReq/phi_stmt_1920/phi_stmt_1920_req
      -- 
    cp_element_group_1242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1240) & cp_elements(1241);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1242), clk => clk, reset => reset); --
    end block;
    phi_stmt_1920_req_13673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1242), ack => phi_stmt_1920_req_2); -- 
    -- CP-element group 1243 merge  place  bypass 
    -- predecessors 1236 1239 1242 
    -- successors 1244 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1919_PhiReqMerge
      -- 
    cp_elements(1243) <= OrReduce(cp_elements(1236) & cp_elements(1239) & cp_elements(1242));
    -- CP-element group 1244 transition  bypass 
    -- predecessors 1243 
    -- successors 1245 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_1919_PhiAck/$entry
      -- 
    cp_elements(1244) <= cp_elements(1243);
    -- CP-element group 1245 transition  place  input  bypass 
    -- predecessors 1244 
    -- successors 228 
    -- members (4) 
      -- 	branch_block_stmt_1659/merge_stmt_1919__exit__
      -- 	branch_block_stmt_1659/assign_stmt_1936_to_assign_stmt_1961__entry__
      -- 	branch_block_stmt_1659/merge_stmt_1919_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_1919_PhiAck/phi_stmt_1920_ack
      -- 
    phi_stmt_1920_ack_13678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1920_ack_0, ack => cp_elements(1245)); -- 
    -- CP-element group 1246 fork  transition  bypass 
    -- predecessors 12 
    -- successors 1247 1251 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/$entry
      -- 
    cp_elements(1246) <= cp_elements(12);
    -- CP-element group 1247 fork  transition  bypass 
    -- predecessors 1246 
    -- successors 1248 1249 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/$entry
      -- 
    cp_elements(1247) <= cp_elements(1246);
    -- CP-element group 1248 transition  bypass 
    -- predecessors 1247 
    -- successors 1250 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/ra
      -- 
    cp_elements(1248) <= cp_elements(1247);
    -- CP-element group 1249 transition  bypass 
    -- predecessors 1247 
    -- successors 1250 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/ca
      -- 
    cp_elements(1249) <= cp_elements(1247);
    -- CP-element group 1250 join  transition  output  bypass 
    -- predecessors 1248 1249 
    -- successors 1263 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_req
      -- 
    cp_element_group_1250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1248) & cp_elements(1249);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1250), clk => clk, reset => reset); --
    end block;
    phi_stmt_2064_req_13728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1250), ack => phi_stmt_2064_req_1); -- 
    -- CP-element group 1251 fork  transition  bypass 
    -- predecessors 1246 
    -- successors 1252 1256 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$entry
      -- 
    cp_elements(1251) <= cp_elements(1246);
    -- CP-element group 1252 fork  transition  bypass 
    -- predecessors 1251 
    -- successors 1253 1254 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$entry
      -- 
    cp_elements(1252) <= cp_elements(1251);
    -- CP-element group 1253 transition  bypass 
    -- predecessors 1252 
    -- successors 1255 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/ra
      -- 
    cp_elements(1253) <= cp_elements(1252);
    -- CP-element group 1254 transition  bypass 
    -- predecessors 1252 
    -- successors 1255 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/ca
      -- 
    cp_elements(1254) <= cp_elements(1252);
    -- CP-element group 1255 join  transition  bypass 
    -- predecessors 1253 1254 
    -- successors 1262 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$exit
      -- 
    cp_element_group_1255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1253) & cp_elements(1254);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1256 fork  transition  bypass 
    -- predecessors 1251 
    -- successors 1257 1259 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/$entry
      -- 
    cp_elements(1256) <= cp_elements(1251);
    -- CP-element group 1257 transition  output  bypass 
    -- predecessors 1256 
    -- successors 1258 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/rr
      -- 
    cp_elements(1257) <= cp_elements(1256);
    rr_13760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1257), ack => type_cast_2063_inst_req_0); -- 
    -- CP-element group 1258 transition  input  bypass 
    -- predecessors 1257 
    -- successors 1261 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/ra
      -- 
    ra_13761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2063_inst_ack_0, ack => cp_elements(1258)); -- 
    -- CP-element group 1259 transition  output  bypass 
    -- predecessors 1256 
    -- successors 1260 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/cr
      -- 
    cp_elements(1259) <= cp_elements(1256);
    cr_13765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1259), ack => type_cast_2063_inst_req_1); -- 
    -- CP-element group 1260 transition  input  bypass 
    -- predecessors 1259 
    -- successors 1261 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/ca
      -- 
    ca_13766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2063_inst_ack_1, ack => cp_elements(1260)); -- 
    -- CP-element group 1261 join  transition  bypass 
    -- predecessors 1258 1260 
    -- successors 1262 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/$exit
      -- 
    cp_element_group_1261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1258) & cp_elements(1260);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1262 join  transition  output  bypass 
    -- predecessors 1255 1261 
    -- successors 1263 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_req
      -- 
    cp_element_group_1262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1255) & cp_elements(1261);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1262), clk => clk, reset => reset); --
    end block;
    phi_stmt_2058_req_13767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1262), ack => phi_stmt_2058_req_1); -- 
    -- CP-element group 1263 join  transition  bypass 
    -- predecessors 1250 1262 
    -- successors 1284 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5x_xpreheader_bbx_xnph7x_xix_xix_xi5_PhiReq/$exit
      -- 
    cp_element_group_1263: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1263"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1250) & cp_elements(1262);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1264 fork  transition  bypass 
    -- predecessors 397 
    -- successors 1265 1271 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/$entry
      -- 
    cp_elements(1264) <= cp_elements(397);
    -- CP-element group 1265 fork  transition  bypass 
    -- predecessors 1264 
    -- successors 1266 1268 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/$entry
      -- 
    cp_elements(1265) <= cp_elements(1264);
    -- CP-element group 1266 transition  output  bypass 
    -- predecessors 1265 
    -- successors 1267 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/rr
      -- 
    cp_elements(1266) <= cp_elements(1265);
    rr_13786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1266), ack => type_cast_2067_inst_req_0); -- 
    -- CP-element group 1267 transition  input  bypass 
    -- predecessors 1266 
    -- successors 1270 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Sample/ra
      -- 
    ra_13787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_0, ack => cp_elements(1267)); -- 
    -- CP-element group 1268 transition  output  bypass 
    -- predecessors 1265 
    -- successors 1269 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/cr
      -- 
    cp_elements(1268) <= cp_elements(1265);
    cr_13791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1268), ack => type_cast_2067_inst_req_1); -- 
    -- CP-element group 1269 transition  input  bypass 
    -- predecessors 1268 
    -- successors 1270 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/Update/ca
      -- 
    ca_13792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_1, ack => cp_elements(1269)); -- 
    -- CP-element group 1270 join  transition  output  bypass 
    -- predecessors 1267 1269 
    -- successors 1283 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_sources/type_cast_2067/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2064/phi_stmt_2064_req
      -- 
    cp_element_group_1270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1267) & cp_elements(1269);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1270), clk => clk, reset => reset); --
    end block;
    phi_stmt_2064_req_13793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1270), ack => phi_stmt_2064_req_0); -- 
    -- CP-element group 1271 fork  transition  bypass 
    -- predecessors 1264 
    -- successors 1272 1278 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$entry
      -- 
    cp_elements(1271) <= cp_elements(1264);
    -- CP-element group 1272 fork  transition  bypass 
    -- predecessors 1271 
    -- successors 1273 1275 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$entry
      -- 
    cp_elements(1272) <= cp_elements(1271);
    -- CP-element group 1273 transition  output  bypass 
    -- predecessors 1272 
    -- successors 1274 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/rr
      -- 
    cp_elements(1273) <= cp_elements(1272);
    rr_13809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1273), ack => type_cast_2061_inst_req_0); -- 
    -- CP-element group 1274 transition  input  bypass 
    -- predecessors 1273 
    -- successors 1277 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Sample/ra
      -- 
    ra_13810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => cp_elements(1274)); -- 
    -- CP-element group 1275 transition  output  bypass 
    -- predecessors 1272 
    -- successors 1276 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/cr
      -- 
    cp_elements(1275) <= cp_elements(1272);
    cr_13814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1275), ack => type_cast_2061_inst_req_1); -- 
    -- CP-element group 1276 transition  input  bypass 
    -- predecessors 1275 
    -- successors 1277 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/Update/ca
      -- 
    ca_13815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => cp_elements(1276)); -- 
    -- CP-element group 1277 join  transition  bypass 
    -- predecessors 1274 1276 
    -- successors 1282 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2061/SplitProtocol/$exit
      -- 
    cp_element_group_1277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1274) & cp_elements(1276);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1278 fork  transition  bypass 
    -- predecessors 1271 
    -- successors 1279 1280 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/$entry
      -- 
    cp_elements(1278) <= cp_elements(1271);
    -- CP-element group 1279 transition  bypass 
    -- predecessors 1278 
    -- successors 1281 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Sample/ra
      -- 
    cp_elements(1279) <= cp_elements(1278);
    -- CP-element group 1280 transition  bypass 
    -- predecessors 1278 
    -- successors 1281 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/Update/ca
      -- 
    cp_elements(1280) <= cp_elements(1278);
    -- CP-element group 1281 join  transition  bypass 
    -- predecessors 1279 1280 
    -- successors 1282 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/type_cast_2063/SplitProtocol/$exit
      -- 
    cp_element_group_1281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1279) & cp_elements(1280);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1282 join  transition  output  bypass 
    -- predecessors 1277 1281 
    -- successors 1283 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/phi_stmt_2058/phi_stmt_2058_req
      -- 
    cp_element_group_1282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1277) & cp_elements(1281);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1282), clk => clk, reset => reset); --
    end block;
    phi_stmt_2058_req_13832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1282), ack => phi_stmt_2058_req_0); -- 
    -- CP-element group 1283 join  transition  bypass 
    -- predecessors 1270 1282 
    -- successors 1284 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_bbx_xnph7x_xix_xix_xi5_PhiReq/$exit
      -- 
    cp_element_group_1283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1270) & cp_elements(1282);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1284 merge  place  bypass 
    -- predecessors 1263 1283 
    -- successors 1285 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2057_PhiReqMerge
      -- 
    cp_elements(1284) <= OrReduce(cp_elements(1263) & cp_elements(1283));
    -- CP-element group 1285 fork  transition  bypass 
    -- predecessors 1284 
    -- successors 1286 1287 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2057_PhiAck/$entry
      -- 
    cp_elements(1285) <= cp_elements(1284);
    -- CP-element group 1286 transition  input  bypass 
    -- predecessors 1285 
    -- successors 1288 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2057_PhiAck/phi_stmt_2058_ack
      -- 
    phi_stmt_2058_ack_13837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2058_ack_0, ack => cp_elements(1286)); -- 
    -- CP-element group 1287 transition  input  bypass 
    -- predecessors 1285 
    -- successors 1288 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2057_PhiAck/phi_stmt_2064_ack
      -- 
    phi_stmt_2064_ack_13838_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2064_ack_0, ack => cp_elements(1287)); -- 
    -- CP-element group 1288 join  transition  bypass 
    -- predecessors 1286 1287 
    -- successors 13 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2057_PhiAck/$exit
      -- 
    cp_element_group_1288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1286) & cp_elements(1287);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1289 fork  transition  bypass 
    -- predecessors 369 
    -- successors 1290 1296 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/$entry
      -- 
    cp_elements(1289) <= cp_elements(369);
    -- CP-element group 1290 fork  transition  bypass 
    -- predecessors 1289 
    -- successors 1291 1293 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$entry
      -- 
    cp_elements(1290) <= cp_elements(1289);
    -- CP-element group 1291 transition  output  bypass 
    -- predecessors 1290 
    -- successors 1292 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/rr
      -- 
    cp_elements(1291) <= cp_elements(1290);
    rr_13869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1291), ack => type_cast_2101_inst_req_0); -- 
    -- CP-element group 1292 transition  input  bypass 
    -- predecessors 1291 
    -- successors 1295 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/ra
      -- 
    ra_13870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_0, ack => cp_elements(1292)); -- 
    -- CP-element group 1293 transition  output  bypass 
    -- predecessors 1290 
    -- successors 1294 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/cr
      -- 
    cp_elements(1293) <= cp_elements(1290);
    cr_13874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1293), ack => type_cast_2101_inst_req_1); -- 
    -- CP-element group 1294 transition  input  bypass 
    -- predecessors 1293 
    -- successors 1295 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/ca
      -- 
    ca_13875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_1, ack => cp_elements(1294)); -- 
    -- CP-element group 1295 join  transition  output  bypass 
    -- predecessors 1292 1294 
    -- successors 1308 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_req
      -- 
    cp_element_group_1295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1292) & cp_elements(1294);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1295), clk => clk, reset => reset); --
    end block;
    phi_stmt_2098_req_13876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1295), ack => phi_stmt_2098_req_0); -- 
    -- CP-element group 1296 fork  transition  bypass 
    -- predecessors 1289 
    -- successors 1297 1303 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/$entry
      -- 
    cp_elements(1296) <= cp_elements(1289);
    -- CP-element group 1297 fork  transition  bypass 
    -- predecessors 1296 
    -- successors 1298 1300 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/$entry
      -- 
    cp_elements(1297) <= cp_elements(1296);
    -- CP-element group 1298 transition  output  bypass 
    -- predecessors 1297 
    -- successors 1299 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/rr
      -- 
    cp_elements(1298) <= cp_elements(1297);
    rr_13892_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1298), ack => type_cast_2095_inst_req_0); -- 
    -- CP-element group 1299 transition  input  bypass 
    -- predecessors 1298 
    -- successors 1302 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/ra
      -- 
    ra_13893_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2095_inst_ack_0, ack => cp_elements(1299)); -- 
    -- CP-element group 1300 transition  output  bypass 
    -- predecessors 1297 
    -- successors 1301 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/cr
      -- 
    cp_elements(1300) <= cp_elements(1297);
    cr_13897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1300), ack => type_cast_2095_inst_req_1); -- 
    -- CP-element group 1301 transition  input  bypass 
    -- predecessors 1300 
    -- successors 1302 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/ca
      -- 
    ca_13898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2095_inst_ack_1, ack => cp_elements(1301)); -- 
    -- CP-element group 1302 join  transition  bypass 
    -- predecessors 1299 1301 
    -- successors 1307 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/$exit
      -- 
    cp_element_group_1302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1299) & cp_elements(1301);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1303 fork  transition  bypass 
    -- predecessors 1296 
    -- successors 1304 1305 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/$entry
      -- 
    cp_elements(1303) <= cp_elements(1296);
    -- CP-element group 1304 transition  bypass 
    -- predecessors 1303 
    -- successors 1306 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/ra
      -- 
    cp_elements(1304) <= cp_elements(1303);
    -- CP-element group 1305 transition  bypass 
    -- predecessors 1303 
    -- successors 1306 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/ca
      -- 
    cp_elements(1305) <= cp_elements(1303);
    -- CP-element group 1306 join  transition  bypass 
    -- predecessors 1304 1305 
    -- successors 1307 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/$exit
      -- 
    cp_element_group_1306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1304) & cp_elements(1305);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1307 join  transition  output  bypass 
    -- predecessors 1302 1306 
    -- successors 1308 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_req
      -- 
    cp_element_group_1307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1302) & cp_elements(1306);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1307), clk => clk, reset => reset); --
    end block;
    phi_stmt_2092_req_13915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1307), ack => phi_stmt_2092_req_0); -- 
    -- CP-element group 1308 join  transition  bypass 
    -- predecessors 1295 1307 
    -- successors 1327 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_bbx_xnphx_xix_xix_xi8_PhiReq/$exit
      -- 
    cp_element_group_1308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1295) & cp_elements(1307);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1309 fork  transition  bypass 
    -- predecessors 14 
    -- successors 1310 1314 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/$entry
      -- 
    cp_elements(1309) <= cp_elements(14);
    -- CP-element group 1310 fork  transition  bypass 
    -- predecessors 1309 
    -- successors 1311 1312 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$entry
      -- 
    cp_elements(1310) <= cp_elements(1309);
    -- CP-element group 1311 transition  bypass 
    -- predecessors 1310 
    -- successors 1313 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/ra
      -- 
    cp_elements(1311) <= cp_elements(1310);
    -- CP-element group 1312 transition  bypass 
    -- predecessors 1310 
    -- successors 1313 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/ca
      -- 
    cp_elements(1312) <= cp_elements(1310);
    -- CP-element group 1313 join  transition  output  bypass 
    -- predecessors 1311 1312 
    -- successors 1326 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2098/phi_stmt_2098_req
      -- 
    cp_element_group_1313: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1313"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1311) & cp_elements(1312);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1313), clk => clk, reset => reset); --
    end block;
    phi_stmt_2098_req_13941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1313), ack => phi_stmt_2098_req_1); -- 
    -- CP-element group 1314 fork  transition  bypass 
    -- predecessors 1309 
    -- successors 1315 1319 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/$entry
      -- 
    cp_elements(1314) <= cp_elements(1309);
    -- CP-element group 1315 fork  transition  bypass 
    -- predecessors 1314 
    -- successors 1316 1317 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/$entry
      -- 
    cp_elements(1315) <= cp_elements(1314);
    -- CP-element group 1316 transition  bypass 
    -- predecessors 1315 
    -- successors 1318 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Sample/ra
      -- 
    cp_elements(1316) <= cp_elements(1315);
    -- CP-element group 1317 transition  bypass 
    -- predecessors 1315 
    -- successors 1318 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/Update/ca
      -- 
    cp_elements(1317) <= cp_elements(1315);
    -- CP-element group 1318 join  transition  bypass 
    -- predecessors 1316 1317 
    -- successors 1325 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2095/SplitProtocol/$exit
      -- 
    cp_element_group_1318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1316) & cp_elements(1317);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1319 fork  transition  bypass 
    -- predecessors 1314 
    -- successors 1320 1322 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/$entry
      -- 
    cp_elements(1319) <= cp_elements(1314);
    -- CP-element group 1320 transition  output  bypass 
    -- predecessors 1319 
    -- successors 1321 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/rr
      -- 
    cp_elements(1320) <= cp_elements(1319);
    rr_13973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1320), ack => type_cast_2097_inst_req_0); -- 
    -- CP-element group 1321 transition  input  bypass 
    -- predecessors 1320 
    -- successors 1324 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Sample/ra
      -- 
    ra_13974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2097_inst_ack_0, ack => cp_elements(1321)); -- 
    -- CP-element group 1322 transition  output  bypass 
    -- predecessors 1319 
    -- successors 1323 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/cr
      -- 
    cp_elements(1322) <= cp_elements(1319);
    cr_13978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1322), ack => type_cast_2097_inst_req_1); -- 
    -- CP-element group 1323 transition  input  bypass 
    -- predecessors 1322 
    -- successors 1324 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/Update/ca
      -- 
    ca_13979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2097_inst_ack_1, ack => cp_elements(1323)); -- 
    -- CP-element group 1324 join  transition  bypass 
    -- predecessors 1321 1323 
    -- successors 1325 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/type_cast_2097/SplitProtocol/$exit
      -- 
    cp_element_group_1324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1321) & cp_elements(1323);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1325 join  transition  output  bypass 
    -- predecessors 1318 1324 
    -- successors 1326 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/phi_stmt_2092/phi_stmt_2092_req
      -- 
    cp_element_group_1325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1318) & cp_elements(1324);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1325), clk => clk, reset => reset); --
    end block;
    phi_stmt_2092_req_13980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1325), ack => phi_stmt_2092_req_1); -- 
    -- CP-element group 1326 join  transition  bypass 
    -- predecessors 1313 1325 
    -- successors 1327 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8x_xpreheader_bbx_xnphx_xix_xix_xi8_PhiReq/$exit
      -- 
    cp_element_group_1326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1313) & cp_elements(1325);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1327 merge  place  bypass 
    -- predecessors 1308 1326 
    -- successors 1328 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2091_PhiReqMerge
      -- 
    cp_elements(1327) <= OrReduce(cp_elements(1308) & cp_elements(1326));
    -- CP-element group 1328 fork  transition  bypass 
    -- predecessors 1327 
    -- successors 1329 1330 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2091_PhiAck/$entry
      -- 
    cp_elements(1328) <= cp_elements(1327);
    -- CP-element group 1329 transition  input  bypass 
    -- predecessors 1328 
    -- successors 1331 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2091_PhiAck/phi_stmt_2092_ack
      -- 
    phi_stmt_2092_ack_13985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2092_ack_0, ack => cp_elements(1329)); -- 
    -- CP-element group 1330 transition  input  bypass 
    -- predecessors 1328 
    -- successors 1331 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2091_PhiAck/phi_stmt_2098_ack
      -- 
    phi_stmt_2098_ack_13986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2098_ack_0, ack => cp_elements(1330)); -- 
    -- CP-element group 1331 join  transition  bypass 
    -- predecessors 1329 1330 
    -- successors 15 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2091_PhiAck/$exit
      -- 
    cp_element_group_1331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1329) & cp_elements(1330);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1332 fork  transition  bypass 
    -- predecessors 371 
    -- successors 1333 1339 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/$entry
      -- 
    cp_elements(1332) <= cp_elements(371);
    -- CP-element group 1333 fork  transition  bypass 
    -- predecessors 1332 
    -- successors 1334 1336 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/$entry
      -- 
    cp_elements(1333) <= cp_elements(1332);
    -- CP-element group 1334 transition  output  bypass 
    -- predecessors 1333 
    -- successors 1335 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Sample/rr
      -- 
    cp_elements(1334) <= cp_elements(1333);
    rr_14009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1334), ack => type_cast_2133_inst_req_0); -- 
    -- CP-element group 1335 transition  input  bypass 
    -- predecessors 1334 
    -- successors 1338 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Sample/ra
      -- 
    ra_14010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_0, ack => cp_elements(1335)); -- 
    -- CP-element group 1336 transition  output  bypass 
    -- predecessors 1333 
    -- successors 1337 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Update/cr
      -- 
    cp_elements(1336) <= cp_elements(1333);
    cr_14014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1336), ack => type_cast_2133_inst_req_1); -- 
    -- CP-element group 1337 transition  input  bypass 
    -- predecessors 1336 
    -- successors 1338 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/Update/ca
      -- 
    ca_14015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_1, ack => cp_elements(1337)); -- 
    -- CP-element group 1338 join  transition  output  bypass 
    -- predecessors 1335 1337 
    -- successors 1345 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_sources/type_cast_2133/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2130/phi_stmt_2130_req
      -- 
    cp_element_group_1338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1335) & cp_elements(1337);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1338), clk => clk, reset => reset); --
    end block;
    phi_stmt_2130_req_14016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1338), ack => phi_stmt_2130_req_0); -- 
    -- CP-element group 1339 fork  transition  bypass 
    -- predecessors 1332 
    -- successors 1340 1342 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$entry
      -- 
    cp_elements(1339) <= cp_elements(1332);
    -- CP-element group 1340 transition  output  bypass 
    -- predecessors 1339 
    -- successors 1341 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/rr
      -- 
    cp_elements(1340) <= cp_elements(1339);
    rr_14032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1340), ack => type_cast_2137_inst_req_0); -- 
    -- CP-element group 1341 transition  input  bypass 
    -- predecessors 1340 
    -- successors 1344 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Sample/ra
      -- 
    ra_14033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2137_inst_ack_0, ack => cp_elements(1341)); -- 
    -- CP-element group 1342 transition  output  bypass 
    -- predecessors 1339 
    -- successors 1343 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/cr
      -- 
    cp_elements(1342) <= cp_elements(1339);
    cr_14037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1342), ack => type_cast_2137_inst_req_1); -- 
    -- CP-element group 1343 transition  input  bypass 
    -- predecessors 1342 
    -- successors 1344 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/Update/ca
      -- 
    ca_14038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2137_inst_ack_1, ack => cp_elements(1343)); -- 
    -- CP-element group 1344 join  transition  output  bypass 
    -- predecessors 1341 1343 
    -- successors 1345 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_sources/type_cast_2137/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/phi_stmt_2134/phi_stmt_2134_req
      -- 
    cp_element_group_1344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1341) & cp_elements(1343);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1344), clk => clk, reset => reset); --
    end block;
    phi_stmt_2134_req_14039_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1344), ack => phi_stmt_2134_req_0); -- 
    -- CP-element group 1345 join  transition  bypass 
    -- predecessors 1338 1344 
    -- successors 1346 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi8_xx_x_crit_edgex_xix_xix_xi11x_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_1345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1338) & cp_elements(1344);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1346 place  bypass 
    -- predecessors 1345 
    -- successors 1347 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2129_PhiReqMerge
      -- 
    cp_elements(1346) <= cp_elements(1345);
    -- CP-element group 1347 fork  transition  bypass 
    -- predecessors 1346 
    -- successors 1348 1349 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2129_PhiAck/$entry
      -- 
    cp_elements(1347) <= cp_elements(1346);
    -- CP-element group 1348 transition  input  bypass 
    -- predecessors 1347 
    -- successors 1350 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2129_PhiAck/phi_stmt_2130_ack
      -- 
    phi_stmt_2130_ack_14044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2130_ack_0, ack => cp_elements(1348)); -- 
    -- CP-element group 1349 transition  input  bypass 
    -- predecessors 1347 
    -- successors 1350 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2129_PhiAck/phi_stmt_2134_ack
      -- 
    phi_stmt_2134_ack_14045_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2134_ack_0, ack => cp_elements(1349)); -- 
    -- CP-element group 1350 join  transition  bypass 
    -- predecessors 1348 1349 
    -- successors 17 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2129_PhiAck/$exit
      -- 
    cp_element_group_1350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1348) & cp_elements(1349);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1351 fork  transition  bypass 
    -- predecessors 349 
    -- successors 1352 1364 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$entry
      -- 
    cp_elements(1351) <= cp_elements(349);
    -- CP-element group 1352 fork  transition  bypass 
    -- predecessors 1351 
    -- successors 1353 1359 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/$entry
      -- 
    cp_elements(1352) <= cp_elements(1351);
    -- CP-element group 1353 fork  transition  bypass 
    -- predecessors 1352 
    -- successors 1354 1356 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/$entry
      -- 
    cp_elements(1353) <= cp_elements(1352);
    -- CP-element group 1354 transition  output  bypass 
    -- predecessors 1353 
    -- successors 1355 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/rr
      -- 
    cp_elements(1354) <= cp_elements(1353);
    rr_14064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1354), ack => type_cast_2144_inst_req_0); -- 
    -- CP-element group 1355 transition  input  bypass 
    -- predecessors 1354 
    -- successors 1358 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/ra
      -- 
    ra_14065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2144_inst_ack_0, ack => cp_elements(1355)); -- 
    -- CP-element group 1356 transition  output  bypass 
    -- predecessors 1353 
    -- successors 1357 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/cr
      -- 
    cp_elements(1356) <= cp_elements(1353);
    cr_14069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1356), ack => type_cast_2144_inst_req_1); -- 
    -- CP-element group 1357 transition  input  bypass 
    -- predecessors 1356 
    -- successors 1358 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/$exit
      -- 
    ca_14070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2144_inst_ack_1, ack => cp_elements(1357)); -- 
    -- CP-element group 1358 join  transition  bypass 
    -- predecessors 1355 1357 
    -- successors 1363 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/$exit
      -- 
    cp_element_group_1358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1355) & cp_elements(1357);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1359 fork  transition  bypass 
    -- predecessors 1352 
    -- successors 1360 1361 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/$entry
      -- 
    cp_elements(1359) <= cp_elements(1352);
    -- CP-element group 1360 transition  bypass 
    -- predecessors 1359 
    -- successors 1362 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1360) <= cp_elements(1359);
    -- CP-element group 1361 transition  bypass 
    -- predecessors 1359 
    -- successors 1362 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/$entry
      -- 
    cp_elements(1361) <= cp_elements(1359);
    -- CP-element group 1362 join  transition  bypass 
    -- predecessors 1360 1361 
    -- successors 1363 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/$exit
      -- 
    cp_element_group_1362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1360) & cp_elements(1361);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1363 join  transition  output  bypass 
    -- predecessors 1358 1362 
    -- successors 1368 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_req
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/$exit
      -- 
    cp_element_group_1363: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1363"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1358) & cp_elements(1362);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1363), clk => clk, reset => reset); --
    end block;
    phi_stmt_2141_req_14087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1363), ack => phi_stmt_2141_req_0); -- 
    -- CP-element group 1364 fork  transition  bypass 
    -- predecessors 1351 
    -- successors 1365 1366 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/$entry
      -- 
    cp_elements(1364) <= cp_elements(1351);
    -- CP-element group 1365 transition  bypass 
    -- predecessors 1364 
    -- successors 1367 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/rr
      -- 
    cp_elements(1365) <= cp_elements(1364);
    -- CP-element group 1366 transition  bypass 
    -- predecessors 1364 
    -- successors 1367 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/$exit
      -- 
    cp_elements(1366) <= cp_elements(1364);
    -- CP-element group 1367 join  transition  output  bypass 
    -- predecessors 1365 1366 
    -- successors 1368 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_req
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/$exit
      -- 
    cp_element_group_1367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1365) & cp_elements(1366);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1367), clk => clk, reset => reset); --
    end block;
    phi_stmt_2147_req_14110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1367), ack => phi_stmt_2147_req_0); -- 
    -- CP-element group 1368 join  transition  bypass 
    -- predecessors 1363 1367 
    -- successors 1389 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi5_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$exit
      -- 
    cp_element_group_1368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1363) & cp_elements(1367);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1369 fork  transition  bypass 
    -- predecessors 17 
    -- successors 1370 1382 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$entry
      -- 
    cp_elements(1369) <= cp_elements(17);
    -- CP-element group 1370 fork  transition  bypass 
    -- predecessors 1369 
    -- successors 1371 1375 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/$entry
      -- 
    cp_elements(1370) <= cp_elements(1369);
    -- CP-element group 1371 fork  transition  bypass 
    -- predecessors 1370 
    -- successors 1372 1373 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/$entry
      -- 
    cp_elements(1371) <= cp_elements(1370);
    -- CP-element group 1372 transition  bypass 
    -- predecessors 1371 
    -- successors 1374 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1372) <= cp_elements(1371);
    -- CP-element group 1373 transition  bypass 
    -- predecessors 1371 
    -- successors 1374 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/Update/$entry
      -- 
    cp_elements(1373) <= cp_elements(1371);
    -- CP-element group 1374 join  transition  bypass 
    -- predecessors 1372 1373 
    -- successors 1381 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2144/$exit
      -- 
    cp_element_group_1374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1372) & cp_elements(1373);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1375 fork  transition  bypass 
    -- predecessors 1370 
    -- successors 1376 1378 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/$entry
      -- 
    cp_elements(1375) <= cp_elements(1370);
    -- CP-element group 1376 transition  output  bypass 
    -- predecessors 1375 
    -- successors 1377 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1376) <= cp_elements(1375);
    rr_14145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1376), ack => type_cast_2146_inst_req_0); -- 
    -- CP-element group 1377 transition  input  bypass 
    -- predecessors 1376 
    -- successors 1380 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Sample/$exit
      -- 
    ra_14146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_0, ack => cp_elements(1377)); -- 
    -- CP-element group 1378 transition  output  bypass 
    -- predecessors 1375 
    -- successors 1379 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/$entry
      -- 
    cp_elements(1378) <= cp_elements(1375);
    cr_14150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1378), ack => type_cast_2146_inst_req_1); -- 
    -- CP-element group 1379 transition  input  bypass 
    -- predecessors 1378 
    -- successors 1380 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/Update/$exit
      -- 
    ca_14151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_1, ack => cp_elements(1379)); -- 
    -- CP-element group 1380 join  transition  bypass 
    -- predecessors 1377 1379 
    -- successors 1381 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/type_cast_2146/$exit
      -- 
    cp_element_group_1380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1377) & cp_elements(1379);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1381 join  transition  output  bypass 
    -- predecessors 1374 1380 
    -- successors 1388 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2141/phi_stmt_2141_req
      -- 
    cp_element_group_1381: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1381"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1374) & cp_elements(1380);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1381), clk => clk, reset => reset); --
    end block;
    phi_stmt_2141_req_14152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1381), ack => phi_stmt_2141_req_1); -- 
    -- CP-element group 1382 fork  transition  bypass 
    -- predecessors 1369 
    -- successors 1383 1385 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/$entry
      -- 
    cp_elements(1382) <= cp_elements(1369);
    -- CP-element group 1383 transition  output  bypass 
    -- predecessors 1382 
    -- successors 1384 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1383) <= cp_elements(1382);
    rr_14168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1383), ack => type_cast_2153_inst_req_0); -- 
    -- CP-element group 1384 transition  input  bypass 
    -- predecessors 1383 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Sample/$exit
      -- 
    ra_14169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2153_inst_ack_0, ack => cp_elements(1384)); -- 
    -- CP-element group 1385 transition  output  bypass 
    -- predecessors 1382 
    -- successors 1386 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/$entry
      -- 
    cp_elements(1385) <= cp_elements(1382);
    cr_14173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1385), ack => type_cast_2153_inst_req_1); -- 
    -- CP-element group 1386 transition  input  bypass 
    -- predecessors 1385 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/Update/$exit
      -- 
    ca_14174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2153_inst_ack_1, ack => cp_elements(1386)); -- 
    -- CP-element group 1387 join  transition  output  bypass 
    -- predecessors 1384 1386 
    -- successors 1388 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_req
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/type_cast_2153/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/phi_stmt_2147_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/phi_stmt_2147/$exit
      -- 
    cp_element_group_1387: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1387"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1384) & cp_elements(1386);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1387), clk => clk, reset => reset); --
    end block;
    phi_stmt_2147_req_14175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1387), ack => phi_stmt_2147_req_1); -- 
    -- CP-element group 1388 join  transition  bypass 
    -- predecessors 1381 1387 
    -- successors 1389 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11x_xloopexit_xx_x_crit_edgex_xix_xix_xi11_PhiReq/$exit
      -- 
    cp_element_group_1388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1381) & cp_elements(1387);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1389 merge  place  bypass 
    -- predecessors 1368 1388 
    -- successors 1390 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2140_PhiReqMerge
      -- 
    cp_elements(1389) <= OrReduce(cp_elements(1368) & cp_elements(1388));
    -- CP-element group 1390 fork  transition  bypass 
    -- predecessors 1389 
    -- successors 1391 1392 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2140_PhiAck/$entry
      -- 
    cp_elements(1390) <= cp_elements(1389);
    -- CP-element group 1391 transition  input  bypass 
    -- predecessors 1390 
    -- successors 1393 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2140_PhiAck/phi_stmt_2141_ack
      -- 
    phi_stmt_2141_ack_14180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2141_ack_0, ack => cp_elements(1391)); -- 
    -- CP-element group 1392 transition  input  bypass 
    -- predecessors 1390 
    -- successors 1393 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2140_PhiAck/phi_stmt_2147_ack
      -- 
    phi_stmt_2147_ack_14181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2147_ack_0, ack => cp_elements(1392)); -- 
    -- CP-element group 1393 join  transition  bypass 
    -- predecessors 1391 1392 
    -- successors 18 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2140_PhiAck/$exit
      -- 
    cp_element_group_1393: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1393"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1391) & cp_elements(1392);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1394 transition  output  bypass 
    -- predecessors 395 
    -- successors 1395 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/rr
      -- 
    cp_elements(1394) <= cp_elements(395);
    rr_14204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1394), ack => type_cast_2180_inst_req_0); -- 
    -- CP-element group 1395 transition  input  bypass 
    -- predecessors 1394 
    -- successors 1398 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/ra
      -- 
    ra_14205_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => cp_elements(1395)); -- 
    -- CP-element group 1396 transition  output  bypass 
    -- predecessors 395 
    -- successors 1397 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/cr
      -- 
    cp_elements(1396) <= cp_elements(395);
    cr_14209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1396), ack => type_cast_2180_inst_req_1); -- 
    -- CP-element group 1397 transition  input  bypass 
    -- predecessors 1396 
    -- successors 1398 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/ca
      -- 
    ca_14210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => cp_elements(1397)); -- 
    -- CP-element group 1398 join  transition  place  output  bypass 
    -- predecessors 1395 1397 
    -- successors 1399 
    -- members (8) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/phi_stmt_2177_req
      -- 	branch_block_stmt_1659/merge_stmt_2176_PhiAck/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/phi_stmt_2177/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi11_xx_xloopexitx_xix_xix_xi13x_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2176_PhiReqMerge
      -- 
    cp_element_group_1398: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1398"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1395) & cp_elements(1397);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1398), clk => clk, reset => reset); --
    end block;
    phi_stmt_2177_req_14211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1398), ack => phi_stmt_2177_req_0); -- 
    -- CP-element group 1399 transition  input  bypass 
    -- predecessors 1398 
    -- successors 20 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2176_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2176_PhiAck/phi_stmt_2177_ack
      -- 
    phi_stmt_2177_ack_14216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2177_ack_0, ack => cp_elements(1399)); -- 
    -- CP-element group 1400 transition  bypass 
    -- predecessors 328 
    -- successors 1402 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/$exit
      -- 
    cp_elements(1400) <= cp_elements(328);
    -- CP-element group 1401 transition  bypass 
    -- predecessors 328 
    -- successors 1402 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/$exit
      -- 
    cp_elements(1401) <= cp_elements(328);
    -- CP-element group 1402 join  transition  output  bypass 
    -- predecessors 1400 1401 
    -- successors 1408 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/$exit
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/$exit
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- 	branch_block_stmt_1659/bb_12_xx_xloopexitx_xix_xix_xi13_PhiReq/$exit
      -- 
    cp_element_group_1402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1400) & cp_elements(1401);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1402), clk => clk, reset => reset); --
    end block;
    phi_stmt_2184_req_14242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1402), ack => phi_stmt_2184_req_0); -- 
    -- CP-element group 1403 transition  output  bypass 
    -- predecessors 20 
    -- successors 1404 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/rr
      -- 
    cp_elements(1403) <= cp_elements(20);
    rr_14261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1403), ack => type_cast_2190_inst_req_0); -- 
    -- CP-element group 1404 transition  input  bypass 
    -- predecessors 1403 
    -- successors 1407 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Sample/ra
      -- 
    ra_14262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_0, ack => cp_elements(1404)); -- 
    -- CP-element group 1405 transition  output  bypass 
    -- predecessors 20 
    -- successors 1406 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/cr
      -- 
    cp_elements(1405) <= cp_elements(20);
    cr_14266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1405), ack => type_cast_2190_inst_req_1); -- 
    -- CP-element group 1406 transition  input  bypass 
    -- predecessors 1405 
    -- successors 1407 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/Update/ca
      -- 
    ca_14267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_1, ack => cp_elements(1406)); -- 
    -- CP-element group 1407 join  transition  output  bypass 
    -- predecessors 1404 1406 
    -- successors 1408 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2190/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13x_xloopexit_xx_xloopexitx_xix_xix_xi13_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- 
    cp_element_group_1407: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1407"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1404) & cp_elements(1406);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1407), clk => clk, reset => reset); --
    end block;
    phi_stmt_2184_req_14268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1407), ack => phi_stmt_2184_req_1); -- 
    -- CP-element group 1408 merge  place  bypass 
    -- predecessors 1402 1407 
    -- successors 1409 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2183_PhiReqMerge
      -- 
    cp_elements(1408) <= OrReduce(cp_elements(1402) & cp_elements(1407));
    -- CP-element group 1409 transition  bypass 
    -- predecessors 1408 
    -- successors 1410 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2183_PhiAck/$entry
      -- 
    cp_elements(1409) <= cp_elements(1408);
    -- CP-element group 1410 fork  transition  place  input  bypass 
    -- predecessors 1409 
    -- successors 1422 1428 
    -- members (7) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16
      -- 	branch_block_stmt_1659/merge_stmt_2183__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2183_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2183_PhiAck/phi_stmt_2184_ack
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- 
    phi_stmt_2184_ack_14273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2184_ack_0, ack => cp_elements(1410)); -- 
    -- CP-element group 1411 fork  transition  bypass 
    -- predecessors 330 
    -- successors 1412 1413 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$entry
      -- 
    cp_elements(1411) <= cp_elements(330);
    -- CP-element group 1412 transition  bypass 
    -- predecessors 1411 
    -- successors 1414 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/ra
      -- 
    cp_elements(1412) <= cp_elements(1411);
    -- CP-element group 1413 transition  bypass 
    -- predecessors 1411 
    -- successors 1414 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/ca
      -- 
    cp_elements(1413) <= cp_elements(1411);
    -- CP-element group 1414 join  transition  bypass 
    -- predecessors 1412 1413 
    -- successors 1421 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$exit
      -- 
    cp_element_group_1414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1412) & cp_elements(1413);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1415 fork  transition  bypass 
    -- predecessors 330 
    -- successors 1416 1418 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$entry
      -- 
    cp_elements(1415) <= cp_elements(330);
    -- CP-element group 1416 transition  output  bypass 
    -- predecessors 1415 
    -- successors 1417 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- 
    cp_elements(1416) <= cp_elements(1415);
    rr_14308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1416), ack => type_cast_2199_inst_req_0); -- 
    -- CP-element group 1417 transition  input  bypass 
    -- predecessors 1416 
    -- successors 1420 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- 
    ra_14309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => cp_elements(1417)); -- 
    -- CP-element group 1418 transition  output  bypass 
    -- predecessors 1415 
    -- successors 1419 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/cr
      -- 
    cp_elements(1418) <= cp_elements(1415);
    cr_14313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1418), ack => type_cast_2199_inst_req_1); -- 
    -- CP-element group 1419 transition  input  bypass 
    -- predecessors 1418 
    -- successors 1420 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/ca
      -- 
    ca_14314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => cp_elements(1419)); -- 
    -- CP-element group 1420 join  transition  bypass 
    -- predecessors 1417 1419 
    -- successors 1421 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$exit
      -- 
    cp_element_group_1420: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1420"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1417) & cp_elements(1419);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1421 join  transition  output  bypass 
    -- predecessors 1414 1420 
    -- successors 1433 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- 	branch_block_stmt_1659/bb_12_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    cp_element_group_1421: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1421"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1414) & cp_elements(1420);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1421), clk => clk, reset => reset); --
    end block;
    phi_stmt_2194_req_14315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1421), ack => phi_stmt_2194_req_1); -- 
    -- CP-element group 1422 fork  transition  bypass 
    -- predecessors 1410 
    -- successors 1423 1425 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$entry
      -- 
    cp_elements(1422) <= cp_elements(1410);
    -- CP-element group 1423 transition  output  bypass 
    -- predecessors 1422 
    -- successors 1424 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/rr
      -- 
    cp_elements(1423) <= cp_elements(1422);
    rr_14334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1423), ack => type_cast_2197_inst_req_0); -- 
    -- CP-element group 1424 transition  input  bypass 
    -- predecessors 1423 
    -- successors 1427 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/ra
      -- 
    ra_14335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_0, ack => cp_elements(1424)); -- 
    -- CP-element group 1425 transition  output  bypass 
    -- predecessors 1422 
    -- successors 1426 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/cr
      -- 
    cp_elements(1425) <= cp_elements(1422);
    cr_14339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1425), ack => type_cast_2197_inst_req_1); -- 
    -- CP-element group 1426 transition  input  bypass 
    -- predecessors 1425 
    -- successors 1427 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/ca
      -- 
    ca_14340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_1, ack => cp_elements(1426)); -- 
    -- CP-element group 1427 join  transition  bypass 
    -- predecessors 1424 1426 
    -- successors 1432 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$exit
      -- 
    cp_element_group_1427: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1427"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1424) & cp_elements(1426);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1428 fork  transition  bypass 
    -- predecessors 1410 
    -- successors 1429 1430 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$entry
      -- 
    cp_elements(1428) <= cp_elements(1410);
    -- CP-element group 1429 transition  bypass 
    -- predecessors 1428 
    -- successors 1431 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- 
    cp_elements(1429) <= cp_elements(1428);
    -- CP-element group 1430 transition  bypass 
    -- predecessors 1428 
    -- successors 1431 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/ca
      -- 
    cp_elements(1430) <= cp_elements(1428);
    -- CP-element group 1431 join  transition  bypass 
    -- predecessors 1429 1430 
    -- successors 1432 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$exit
      -- 
    cp_element_group_1431: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1431"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1429) & cp_elements(1430);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1432 join  transition  output  bypass 
    -- predecessors 1427 1431 
    -- successors 1433 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi13_udiv32x_xexitx_xpreheaderx_xix_xi16_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    cp_element_group_1432: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1432"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1427) & cp_elements(1431);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1432), clk => clk, reset => reset); --
    end block;
    phi_stmt_2194_req_14357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1432), ack => phi_stmt_2194_req_0); -- 
    -- CP-element group 1433 merge  place  bypass 
    -- predecessors 1421 1432 
    -- successors 1434 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2193_PhiReqMerge
      -- 
    cp_elements(1433) <= OrReduce(cp_elements(1421) & cp_elements(1432));
    -- CP-element group 1434 transition  bypass 
    -- predecessors 1433 
    -- successors 1435 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2193_PhiAck/$entry
      -- 
    cp_elements(1434) <= cp_elements(1433);
    -- CP-element group 1435 transition  place  input  bypass 
    -- predecessors 1434 
    -- successors 398 
    -- members (4) 
      -- 	branch_block_stmt_1659/merge_stmt_2193__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2206_to_assign_stmt_2225__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2193_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2193_PhiAck/phi_stmt_2194_ack
      -- 
    phi_stmt_2194_ack_14362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2194_ack_0, ack => cp_elements(1435)); -- 
    -- CP-element group 1436 fork  transition  bypass 
    -- predecessors 454 
    -- successors 1437 1443 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/$entry
      -- 
    cp_elements(1436) <= cp_elements(454);
    -- CP-element group 1437 fork  transition  bypass 
    -- predecessors 1436 
    -- successors 1438 1440 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/$entry
      -- 
    cp_elements(1437) <= cp_elements(1436);
    -- CP-element group 1438 transition  output  bypass 
    -- predecessors 1437 
    -- successors 1439 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/rr
      -- 
    cp_elements(1438) <= cp_elements(1437);
    rr_14393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1438), ack => type_cast_2238_inst_req_0); -- 
    -- CP-element group 1439 transition  input  bypass 
    -- predecessors 1438 
    -- successors 1442 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/ra
      -- 
    ra_14394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_0, ack => cp_elements(1439)); -- 
    -- CP-element group 1440 transition  output  bypass 
    -- predecessors 1437 
    -- successors 1441 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/cr
      -- 
    cp_elements(1440) <= cp_elements(1437);
    cr_14398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1440), ack => type_cast_2238_inst_req_1); -- 
    -- CP-element group 1441 transition  input  bypass 
    -- predecessors 1440 
    -- successors 1442 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/ca
      -- 
    ca_14399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_1, ack => cp_elements(1441)); -- 
    -- CP-element group 1442 join  transition  output  bypass 
    -- predecessors 1439 1441 
    -- successors 1455 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_req
      -- 
    cp_element_group_1442: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1442"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1439) & cp_elements(1441);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1442), clk => clk, reset => reset); --
    end block;
    phi_stmt_2235_req_14400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1442), ack => phi_stmt_2235_req_0); -- 
    -- CP-element group 1443 fork  transition  bypass 
    -- predecessors 1436 
    -- successors 1444 1450 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/$entry
      -- 
    cp_elements(1443) <= cp_elements(1436);
    -- CP-element group 1444 fork  transition  bypass 
    -- predecessors 1443 
    -- successors 1445 1447 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/$entry
      -- 
    cp_elements(1444) <= cp_elements(1443);
    -- CP-element group 1445 transition  output  bypass 
    -- predecessors 1444 
    -- successors 1446 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/rr
      -- 
    cp_elements(1445) <= cp_elements(1444);
    rr_14416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1445), ack => type_cast_2245_inst_req_0); -- 
    -- CP-element group 1446 transition  input  bypass 
    -- predecessors 1445 
    -- successors 1449 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/ra
      -- 
    ra_14417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2245_inst_ack_0, ack => cp_elements(1446)); -- 
    -- CP-element group 1447 transition  output  bypass 
    -- predecessors 1444 
    -- successors 1448 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/cr
      -- 
    cp_elements(1447) <= cp_elements(1444);
    cr_14421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1447), ack => type_cast_2245_inst_req_1); -- 
    -- CP-element group 1448 transition  input  bypass 
    -- predecessors 1447 
    -- successors 1449 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/ca
      -- 
    ca_14422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2245_inst_ack_1, ack => cp_elements(1448)); -- 
    -- CP-element group 1449 join  transition  bypass 
    -- predecessors 1446 1448 
    -- successors 1454 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/$exit
      -- 
    cp_element_group_1449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1446) & cp_elements(1448);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1450 fork  transition  bypass 
    -- predecessors 1443 
    -- successors 1451 1452 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/$entry
      -- 
    cp_elements(1450) <= cp_elements(1443);
    -- CP-element group 1451 transition  bypass 
    -- predecessors 1450 
    -- successors 1453 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/ra
      -- 
    cp_elements(1451) <= cp_elements(1450);
    -- CP-element group 1452 transition  bypass 
    -- predecessors 1450 
    -- successors 1453 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/ca
      -- 
    cp_elements(1452) <= cp_elements(1450);
    -- CP-element group 1453 join  transition  bypass 
    -- predecessors 1451 1452 
    -- successors 1454 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/$exit
      -- 
    cp_element_group_1453: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1453"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1451) & cp_elements(1452);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1454 join  transition  output  bypass 
    -- predecessors 1449 1453 
    -- successors 1455 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_req
      -- 
    cp_element_group_1454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1449) & cp_elements(1453);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1454), clk => clk, reset => reset); --
    end block;
    phi_stmt_2242_req_14439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1454), ack => phi_stmt_2242_req_0); -- 
    -- CP-element group 1455 join  transition  bypass 
    -- predecessors 1442 1454 
    -- successors 1474 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xix_xi20_PhiReq/$exit
      -- 
    cp_element_group_1455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1442) & cp_elements(1454);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1456 fork  transition  bypass 
    -- predecessors 21 
    -- successors 1457 1461 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/$entry
      -- 
    cp_elements(1456) <= cp_elements(21);
    -- CP-element group 1457 fork  transition  bypass 
    -- predecessors 1456 
    -- successors 1458 1459 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/$entry
      -- 
    cp_elements(1457) <= cp_elements(1456);
    -- CP-element group 1458 transition  bypass 
    -- predecessors 1457 
    -- successors 1460 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Sample/ra
      -- 
    cp_elements(1458) <= cp_elements(1457);
    -- CP-element group 1459 transition  bypass 
    -- predecessors 1457 
    -- successors 1460 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/Update/ca
      -- 
    cp_elements(1459) <= cp_elements(1457);
    -- CP-element group 1460 join  transition  output  bypass 
    -- predecessors 1458 1459 
    -- successors 1473 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_sources/type_cast_2238/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2235/phi_stmt_2235_req
      -- 
    cp_element_group_1460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1458) & cp_elements(1459);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1460), clk => clk, reset => reset); --
    end block;
    phi_stmt_2235_req_14465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1460), ack => phi_stmt_2235_req_1); -- 
    -- CP-element group 1461 fork  transition  bypass 
    -- predecessors 1456 
    -- successors 1462 1466 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/$entry
      -- 
    cp_elements(1461) <= cp_elements(1456);
    -- CP-element group 1462 fork  transition  bypass 
    -- predecessors 1461 
    -- successors 1463 1464 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/$entry
      -- 
    cp_elements(1462) <= cp_elements(1461);
    -- CP-element group 1463 transition  bypass 
    -- predecessors 1462 
    -- successors 1465 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Sample/ra
      -- 
    cp_elements(1463) <= cp_elements(1462);
    -- CP-element group 1464 transition  bypass 
    -- predecessors 1462 
    -- successors 1465 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/Update/ca
      -- 
    cp_elements(1464) <= cp_elements(1462);
    -- CP-element group 1465 join  transition  bypass 
    -- predecessors 1463 1464 
    -- successors 1472 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2245/SplitProtocol/$exit
      -- 
    cp_element_group_1465: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1465"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1463) & cp_elements(1464);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1465), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1466 fork  transition  bypass 
    -- predecessors 1461 
    -- successors 1467 1469 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/$entry
      -- 
    cp_elements(1466) <= cp_elements(1461);
    -- CP-element group 1467 transition  output  bypass 
    -- predecessors 1466 
    -- successors 1468 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/rr
      -- 
    cp_elements(1467) <= cp_elements(1466);
    rr_14497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1467), ack => type_cast_2247_inst_req_0); -- 
    -- CP-element group 1468 transition  input  bypass 
    -- predecessors 1467 
    -- successors 1471 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Sample/ra
      -- 
    ra_14498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_0, ack => cp_elements(1468)); -- 
    -- CP-element group 1469 transition  output  bypass 
    -- predecessors 1466 
    -- successors 1470 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/cr
      -- 
    cp_elements(1469) <= cp_elements(1466);
    cr_14502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1469), ack => type_cast_2247_inst_req_1); -- 
    -- CP-element group 1470 transition  input  bypass 
    -- predecessors 1469 
    -- successors 1471 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/Update/ca
      -- 
    ca_14503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_1, ack => cp_elements(1470)); -- 
    -- CP-element group 1471 join  transition  bypass 
    -- predecessors 1468 1470 
    -- successors 1472 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/type_cast_2247/SplitProtocol/$exit
      -- 
    cp_element_group_1471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1468) & cp_elements(1470);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1472 join  transition  output  bypass 
    -- predecessors 1465 1471 
    -- successors 1473 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/phi_stmt_2242/phi_stmt_2242_req
      -- 
    cp_element_group_1472: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1472"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1465) & cp_elements(1471);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1472), clk => clk, reset => reset); --
    end block;
    phi_stmt_2242_req_14504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1472), ack => phi_stmt_2242_req_1); -- 
    -- CP-element group 1473 join  transition  bypass 
    -- predecessors 1460 1472 
    -- successors 1474 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20x_xpreheader_udiv32x_xexitx_xix_xi20_PhiReq/$exit
      -- 
    cp_element_group_1473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1460) & cp_elements(1472);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1474 merge  place  bypass 
    -- predecessors 1455 1473 
    -- successors 1475 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2234_PhiReqMerge
      -- 
    cp_elements(1474) <= OrReduce(cp_elements(1455) & cp_elements(1473));
    -- CP-element group 1475 fork  transition  bypass 
    -- predecessors 1474 
    -- successors 1476 1477 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2234_PhiAck/$entry
      -- 
    cp_elements(1475) <= cp_elements(1474);
    -- CP-element group 1476 transition  input  bypass 
    -- predecessors 1475 
    -- successors 1478 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2234_PhiAck/phi_stmt_2235_ack
      -- 
    phi_stmt_2235_ack_14509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2235_ack_0, ack => cp_elements(1476)); -- 
    -- CP-element group 1477 transition  input  bypass 
    -- predecessors 1475 
    -- successors 1478 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2234_PhiAck/phi_stmt_2242_ack
      -- 
    phi_stmt_2242_ack_14510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2242_ack_0, ack => cp_elements(1477)); -- 
    -- CP-element group 1478 join  transition  bypass 
    -- predecessors 1476 1477 
    -- successors 22 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2234_PhiAck/$exit
      -- 
    cp_element_group_1478: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1478"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1476) & cp_elements(1477);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1478), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1479 fork  transition  bypass 
    -- predecessors 456 
    -- successors 1480 1486 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/$entry
      -- 
    cp_elements(1479) <= cp_elements(456);
    -- CP-element group 1480 fork  transition  bypass 
    -- predecessors 1479 
    -- successors 1481 1483 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/$entry
      -- 
    cp_elements(1480) <= cp_elements(1479);
    -- CP-element group 1481 transition  output  bypass 
    -- predecessors 1480 
    -- successors 1482 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Sample/rr
      -- 
    cp_elements(1481) <= cp_elements(1480);
    rr_14533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1481), ack => type_cast_2296_inst_req_0); -- 
    -- CP-element group 1482 transition  input  bypass 
    -- predecessors 1481 
    -- successors 1485 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Sample/ra
      -- 
    ra_14534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2296_inst_ack_0, ack => cp_elements(1482)); -- 
    -- CP-element group 1483 transition  output  bypass 
    -- predecessors 1480 
    -- successors 1484 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Update/cr
      -- 
    cp_elements(1483) <= cp_elements(1480);
    cr_14538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1483), ack => type_cast_2296_inst_req_1); -- 
    -- CP-element group 1484 transition  input  bypass 
    -- predecessors 1483 
    -- successors 1485 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/Update/ca
      -- 
    ca_14539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2296_inst_ack_1, ack => cp_elements(1484)); -- 
    -- CP-element group 1485 join  transition  output  bypass 
    -- predecessors 1482 1484 
    -- successors 1492 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_sources/type_cast_2296/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2293/phi_stmt_2293_req
      -- 
    cp_element_group_1485: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1485"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1482) & cp_elements(1484);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1485), clk => clk, reset => reset); --
    end block;
    phi_stmt_2293_req_14540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1485), ack => phi_stmt_2293_req_0); -- 
    -- CP-element group 1486 fork  transition  bypass 
    -- predecessors 1479 
    -- successors 1487 1489 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/$entry
      -- 
    cp_elements(1486) <= cp_elements(1479);
    -- CP-element group 1487 transition  output  bypass 
    -- predecessors 1486 
    -- successors 1488 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/rr
      -- 
    cp_elements(1487) <= cp_elements(1486);
    rr_14556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1487), ack => type_cast_2300_inst_req_0); -- 
    -- CP-element group 1488 transition  input  bypass 
    -- predecessors 1487 
    -- successors 1491 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Sample/ra
      -- 
    ra_14557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_0, ack => cp_elements(1488)); -- 
    -- CP-element group 1489 transition  output  bypass 
    -- predecessors 1486 
    -- successors 1490 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/cr
      -- 
    cp_elements(1489) <= cp_elements(1486);
    cr_14561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1489), ack => type_cast_2300_inst_req_1); -- 
    -- CP-element group 1490 transition  input  bypass 
    -- predecessors 1489 
    -- successors 1491 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/Update/ca
      -- 
    ca_14562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_1, ack => cp_elements(1490)); -- 
    -- CP-element group 1491 join  transition  output  bypass 
    -- predecessors 1488 1490 
    -- successors 1492 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_sources/type_cast_2300/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/phi_stmt_2297/phi_stmt_2297_req
      -- 
    cp_element_group_1491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1488) & cp_elements(1490);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1491), clk => clk, reset => reset); --
    end block;
    phi_stmt_2297_req_14563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1491), ack => phi_stmt_2297_req_0); -- 
    -- CP-element group 1492 join  transition  bypass 
    -- predecessors 1485 1491 
    -- successors 1493 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi20_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_PhiReq/$exit
      -- 
    cp_element_group_1492: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1492"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1485) & cp_elements(1491);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1492), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1493 place  bypass 
    -- predecessors 1492 
    -- successors 1494 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2292_PhiReqMerge
      -- 
    cp_elements(1493) <= cp_elements(1492);
    -- CP-element group 1494 fork  transition  bypass 
    -- predecessors 1493 
    -- successors 1495 1496 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2292_PhiAck/$entry
      -- 
    cp_elements(1494) <= cp_elements(1493);
    -- CP-element group 1495 transition  input  bypass 
    -- predecessors 1494 
    -- successors 1497 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2292_PhiAck/phi_stmt_2293_ack
      -- 
    phi_stmt_2293_ack_14568_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2293_ack_0, ack => cp_elements(1495)); -- 
    -- CP-element group 1496 transition  input  bypass 
    -- predecessors 1494 
    -- successors 1497 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2292_PhiAck/phi_stmt_2297_ack
      -- 
    phi_stmt_2297_ack_14569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2297_ack_0, ack => cp_elements(1496)); -- 
    -- CP-element group 1497 join  transition  bypass 
    -- predecessors 1495 1496 
    -- successors 24 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2292_PhiAck/$exit
      -- 
    cp_element_group_1497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1495) & cp_elements(1496);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1498 fork  transition  bypass 
    -- predecessors 422 
    -- successors 1499 1511 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/$entry
      -- 
    cp_elements(1498) <= cp_elements(422);
    -- CP-element group 1499 fork  transition  bypass 
    -- predecessors 1498 
    -- successors 1500 1504 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/$entry
      -- 
    cp_elements(1499) <= cp_elements(1498);
    -- CP-element group 1500 fork  transition  bypass 
    -- predecessors 1499 
    -- successors 1501 1502 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/$entry
      -- 
    cp_elements(1500) <= cp_elements(1499);
    -- CP-element group 1501 transition  bypass 
    -- predecessors 1500 
    -- successors 1503 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/ra
      -- 
    cp_elements(1501) <= cp_elements(1500);
    -- CP-element group 1502 transition  bypass 
    -- predecessors 1500 
    -- successors 1503 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/ca
      -- 
    cp_elements(1502) <= cp_elements(1500);
    -- CP-element group 1503 join  transition  bypass 
    -- predecessors 1501 1502 
    -- successors 1510 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/$exit
      -- 
    cp_element_group_1503: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1503"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1501) & cp_elements(1502);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1504 fork  transition  bypass 
    -- predecessors 1499 
    -- successors 1505 1507 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/$entry
      -- 
    cp_elements(1504) <= cp_elements(1499);
    -- CP-element group 1505 transition  output  bypass 
    -- predecessors 1504 
    -- successors 1506 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/rr
      -- 
    cp_elements(1505) <= cp_elements(1504);
    rr_14604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1505), ack => type_cast_2331_inst_req_0); -- 
    -- CP-element group 1506 transition  input  bypass 
    -- predecessors 1505 
    -- successors 1509 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/ra
      -- 
    ra_14605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_0, ack => cp_elements(1506)); -- 
    -- CP-element group 1507 transition  output  bypass 
    -- predecessors 1504 
    -- successors 1508 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/cr
      -- 
    cp_elements(1507) <= cp_elements(1504);
    cr_14609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1507), ack => type_cast_2331_inst_req_1); -- 
    -- CP-element group 1508 transition  input  bypass 
    -- predecessors 1507 
    -- successors 1509 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/ca
      -- 
    ca_14610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_1, ack => cp_elements(1508)); -- 
    -- CP-element group 1509 join  transition  bypass 
    -- predecessors 1506 1508 
    -- successors 1510 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/$exit
      -- 
    cp_element_group_1509: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1509"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1506) & cp_elements(1508);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1509), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1510 join  transition  output  bypass 
    -- predecessors 1503 1509 
    -- successors 1523 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_req
      -- 
    cp_element_group_1510: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1510"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1503) & cp_elements(1509);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1510), clk => clk, reset => reset); --
    end block;
    phi_stmt_2326_req_14611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1510), ack => phi_stmt_2326_req_1); -- 
    -- CP-element group 1511 fork  transition  bypass 
    -- predecessors 1498 
    -- successors 1512 1516 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/$entry
      -- 
    cp_elements(1511) <= cp_elements(1498);
    -- CP-element group 1512 fork  transition  bypass 
    -- predecessors 1511 
    -- successors 1513 1514 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/$entry
      -- 
    cp_elements(1512) <= cp_elements(1511);
    -- CP-element group 1513 transition  bypass 
    -- predecessors 1512 
    -- successors 1515 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/ra
      -- 
    cp_elements(1513) <= cp_elements(1512);
    -- CP-element group 1514 transition  bypass 
    -- predecessors 1512 
    -- successors 1515 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/ca
      -- 
    cp_elements(1514) <= cp_elements(1512);
    -- CP-element group 1515 join  transition  bypass 
    -- predecessors 1513 1514 
    -- successors 1522 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/$exit
      -- 
    cp_element_group_1515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1513) & cp_elements(1514);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1516 fork  transition  bypass 
    -- predecessors 1511 
    -- successors 1517 1519 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/$entry
      -- 
    cp_elements(1516) <= cp_elements(1511);
    -- CP-element group 1517 transition  output  bypass 
    -- predecessors 1516 
    -- successors 1518 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/rr
      -- 
    cp_elements(1517) <= cp_elements(1516);
    rr_14643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1517), ack => type_cast_2337_inst_req_0); -- 
    -- CP-element group 1518 transition  input  bypass 
    -- predecessors 1517 
    -- successors 1521 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/ra
      -- 
    ra_14644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2337_inst_ack_0, ack => cp_elements(1518)); -- 
    -- CP-element group 1519 transition  output  bypass 
    -- predecessors 1516 
    -- successors 1520 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/cr
      -- 
    cp_elements(1519) <= cp_elements(1516);
    cr_14648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1519), ack => type_cast_2337_inst_req_1); -- 
    -- CP-element group 1520 transition  input  bypass 
    -- predecessors 1519 
    -- successors 1521 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/ca
      -- 
    ca_14649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2337_inst_ack_1, ack => cp_elements(1520)); -- 
    -- CP-element group 1521 join  transition  bypass 
    -- predecessors 1518 1520 
    -- successors 1522 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/$exit
      -- 
    cp_element_group_1521: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1521"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1518) & cp_elements(1520);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1521), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1522 join  transition  output  bypass 
    -- predecessors 1515 1521 
    -- successors 1523 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_req
      -- 
    cp_element_group_1522: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1522"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1515) & cp_elements(1521);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1522), clk => clk, reset => reset); --
    end block;
    phi_stmt_2332_req_14650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1522), ack => phi_stmt_2332_req_1); -- 
    -- CP-element group 1523 join  transition  bypass 
    -- predecessors 1510 1522 
    -- successors 1550 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi16_xx_xcritedgex_xix_xi29_PhiReq/$exit
      -- 
    cp_element_group_1523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1510) & cp_elements(1522);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1524 fork  transition  bypass 
    -- predecessors 474 
    -- successors 1525 1537 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/$entry
      -- 
    cp_elements(1524) <= cp_elements(474);
    -- CP-element group 1525 fork  transition  bypass 
    -- predecessors 1524 
    -- successors 1526 1532 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/$entry
      -- 
    cp_elements(1525) <= cp_elements(1524);
    -- CP-element group 1526 fork  transition  bypass 
    -- predecessors 1525 
    -- successors 1527 1529 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/$entry
      -- 
    cp_elements(1526) <= cp_elements(1525);
    -- CP-element group 1527 transition  output  bypass 
    -- predecessors 1526 
    -- successors 1528 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/rr
      -- 
    cp_elements(1527) <= cp_elements(1526);
    rr_14669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1527), ack => type_cast_2329_inst_req_0); -- 
    -- CP-element group 1528 transition  input  bypass 
    -- predecessors 1527 
    -- successors 1531 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Sample/ra
      -- 
    ra_14670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2329_inst_ack_0, ack => cp_elements(1528)); -- 
    -- CP-element group 1529 transition  output  bypass 
    -- predecessors 1526 
    -- successors 1530 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/cr
      -- 
    cp_elements(1529) <= cp_elements(1526);
    cr_14674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1529), ack => type_cast_2329_inst_req_1); -- 
    -- CP-element group 1530 transition  input  bypass 
    -- predecessors 1529 
    -- successors 1531 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/Update/ca
      -- 
    ca_14675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2329_inst_ack_1, ack => cp_elements(1530)); -- 
    -- CP-element group 1531 join  transition  bypass 
    -- predecessors 1528 1530 
    -- successors 1536 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2329/SplitProtocol/$exit
      -- 
    cp_element_group_1531: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1531"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1528) & cp_elements(1530);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1531), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1532 fork  transition  bypass 
    -- predecessors 1525 
    -- successors 1533 1534 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/$entry
      -- 
    cp_elements(1532) <= cp_elements(1525);
    -- CP-element group 1533 transition  bypass 
    -- predecessors 1532 
    -- successors 1535 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Sample/ra
      -- 
    cp_elements(1533) <= cp_elements(1532);
    -- CP-element group 1534 transition  bypass 
    -- predecessors 1532 
    -- successors 1535 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/Update/ca
      -- 
    cp_elements(1534) <= cp_elements(1532);
    -- CP-element group 1535 join  transition  bypass 
    -- predecessors 1533 1534 
    -- successors 1536 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/type_cast_2331/SplitProtocol/$exit
      -- 
    cp_element_group_1535: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1535"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1533) & cp_elements(1534);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1535), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1536 join  transition  output  bypass 
    -- predecessors 1531 1535 
    -- successors 1549 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2326/phi_stmt_2326_req
      -- 
    cp_element_group_1536: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1536"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1531) & cp_elements(1535);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1536), clk => clk, reset => reset); --
    end block;
    phi_stmt_2326_req_14692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1536), ack => phi_stmt_2326_req_0); -- 
    -- CP-element group 1537 fork  transition  bypass 
    -- predecessors 1524 
    -- successors 1538 1544 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/$entry
      -- 
    cp_elements(1537) <= cp_elements(1524);
    -- CP-element group 1538 fork  transition  bypass 
    -- predecessors 1537 
    -- successors 1539 1541 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/$entry
      -- 
    cp_elements(1538) <= cp_elements(1537);
    -- CP-element group 1539 transition  output  bypass 
    -- predecessors 1538 
    -- successors 1540 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/rr
      -- 
    cp_elements(1539) <= cp_elements(1538);
    rr_14708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1539), ack => type_cast_2335_inst_req_0); -- 
    -- CP-element group 1540 transition  input  bypass 
    -- predecessors 1539 
    -- successors 1543 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Sample/ra
      -- 
    ra_14709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_0, ack => cp_elements(1540)); -- 
    -- CP-element group 1541 transition  output  bypass 
    -- predecessors 1538 
    -- successors 1542 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/cr
      -- 
    cp_elements(1541) <= cp_elements(1538);
    cr_14713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1541), ack => type_cast_2335_inst_req_1); -- 
    -- CP-element group 1542 transition  input  bypass 
    -- predecessors 1541 
    -- successors 1543 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/Update/ca
      -- 
    ca_14714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_1, ack => cp_elements(1542)); -- 
    -- CP-element group 1543 join  transition  bypass 
    -- predecessors 1540 1542 
    -- successors 1548 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2335/SplitProtocol/$exit
      -- 
    cp_element_group_1543: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1543"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1540) & cp_elements(1542);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1543), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1544 fork  transition  bypass 
    -- predecessors 1537 
    -- successors 1545 1546 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/$entry
      -- 
    cp_elements(1544) <= cp_elements(1537);
    -- CP-element group 1545 transition  bypass 
    -- predecessors 1544 
    -- successors 1547 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Sample/ra
      -- 
    cp_elements(1545) <= cp_elements(1544);
    -- CP-element group 1546 transition  bypass 
    -- predecessors 1544 
    -- successors 1547 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/Update/ca
      -- 
    cp_elements(1546) <= cp_elements(1544);
    -- CP-element group 1547 join  transition  bypass 
    -- predecessors 1545 1546 
    -- successors 1548 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/type_cast_2337/SplitProtocol/$exit
      -- 
    cp_element_group_1547: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1547"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1545) & cp_elements(1546);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1547), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1548 join  transition  output  bypass 
    -- predecessors 1543 1547 
    -- successors 1549 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/phi_stmt_2332/phi_stmt_2332_req
      -- 
    cp_element_group_1548: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1548"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1543) & cp_elements(1547);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1548), clk => clk, reset => reset); --
    end block;
    phi_stmt_2332_req_14731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1548), ack => phi_stmt_2332_req_0); -- 
    -- CP-element group 1549 join  transition  bypass 
    -- predecessors 1536 1548 
    -- successors 1550 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi25_xx_xcritedgex_xix_xi29_PhiReq/$exit
      -- 
    cp_element_group_1549: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1549"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1536) & cp_elements(1548);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1549), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1550 merge  place  bypass 
    -- predecessors 1523 1549 
    -- successors 1551 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2325_PhiReqMerge
      -- 
    cp_elements(1550) <= OrReduce(cp_elements(1523) & cp_elements(1549));
    -- CP-element group 1551 fork  transition  bypass 
    -- predecessors 1550 
    -- successors 1552 1553 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2325_PhiAck/$entry
      -- 
    cp_elements(1551) <= cp_elements(1550);
    -- CP-element group 1552 transition  input  bypass 
    -- predecessors 1551 
    -- successors 1554 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2325_PhiAck/phi_stmt_2326_ack
      -- 
    phi_stmt_2326_ack_14736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2326_ack_0, ack => cp_elements(1552)); -- 
    -- CP-element group 1553 transition  input  bypass 
    -- predecessors 1551 
    -- successors 1554 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2325_PhiAck/phi_stmt_2332_ack
      -- 
    phi_stmt_2332_ack_14737_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2332_ack_0, ack => cp_elements(1553)); -- 
    -- CP-element group 1554 join  transition  bypass 
    -- predecessors 1552 1553 
    -- successors 25 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2325_PhiAck/$exit
      -- 
    cp_element_group_1554: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1554"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1552) & cp_elements(1553);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1554), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1555 transition  bypass 
    -- predecessors 258 
    -- successors 1557 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/ra
      -- 
    cp_elements(1555) <= cp_elements(258);
    -- CP-element group 1556 transition  bypass 
    -- predecessors 258 
    -- successors 1557 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/ca
      -- 
    cp_elements(1556) <= cp_elements(258);
    -- CP-element group 1557 join  transition  output  bypass 
    -- predecessors 1555 1556 
    -- successors 1563 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_11_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_req
      -- 
    cp_element_group_1557: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1557"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1555) & cp_elements(1556);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1557), clk => clk, reset => reset); --
    end block;
    phi_stmt_2373_req_14763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1557), ack => phi_stmt_2373_req_1); -- 
    -- CP-element group 1558 transition  output  bypass 
    -- predecessors 498 
    -- successors 1559 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/rr
      -- 
    cp_elements(1558) <= cp_elements(498);
    rr_14782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1558), ack => type_cast_2376_inst_req_0); -- 
    -- CP-element group 1559 transition  input  bypass 
    -- predecessors 1558 
    -- successors 1562 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Sample/ra
      -- 
    ra_14783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_0, ack => cp_elements(1559)); -- 
    -- CP-element group 1560 transition  output  bypass 
    -- predecessors 498 
    -- successors 1561 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/cr
      -- 
    cp_elements(1560) <= cp_elements(498);
    cr_14787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1560), ack => type_cast_2376_inst_req_1); -- 
    -- CP-element group 1561 transition  input  bypass 
    -- predecessors 1560 
    -- successors 1562 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/Update/ca
      -- 
    ca_14788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_1, ack => cp_elements(1561)); -- 
    -- CP-element group 1562 join  transition  output  bypass 
    -- predecessors 1559 1561 
    -- successors 1563 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_sources/type_cast_2376/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi29_omega_calcx_xexit_PhiReq/phi_stmt_2373/phi_stmt_2373_req
      -- 
    cp_element_group_1562: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1562"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1559) & cp_elements(1561);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1562), clk => clk, reset => reset); --
    end block;
    phi_stmt_2373_req_14789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1562), ack => phi_stmt_2373_req_0); -- 
    -- CP-element group 1563 merge  place  bypass 
    -- predecessors 1557 1562 
    -- successors 1564 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2372_PhiReqMerge
      -- 
    cp_elements(1563) <= OrReduce(cp_elements(1557) & cp_elements(1562));
    -- CP-element group 1564 transition  bypass 
    -- predecessors 1563 
    -- successors 1565 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2372_PhiAck/$entry
      -- 
    cp_elements(1564) <= cp_elements(1563);
    -- CP-element group 1565 transition  place  input  bypass 
    -- predecessors 1564 
    -- successors 499 
    -- members (4) 
      -- 	branch_block_stmt_1659/merge_stmt_2372__exit__
      -- 	branch_block_stmt_1659/assign_stmt_2385_to_assign_stmt_2406__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2372_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2372_PhiAck/phi_stmt_2373_ack
      -- 
    phi_stmt_2373_ack_14794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2373_ack_0, ack => cp_elements(1565)); -- 
    -- CP-element group 1566 fork  transition  bypass 
    -- predecessors 29 
    -- successors 1567 1579 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1566) <= cp_elements(29);
    -- CP-element group 1567 fork  transition  bypass 
    -- predecessors 1566 
    -- successors 1568 1572 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- 
    cp_elements(1567) <= cp_elements(1566);
    -- CP-element group 1568 fork  transition  bypass 
    -- predecessors 1567 
    -- successors 1569 1570 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$entry
      -- 
    cp_elements(1568) <= cp_elements(1567);
    -- CP-element group 1569 transition  bypass 
    -- predecessors 1568 
    -- successors 1571 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/ra
      -- 
    cp_elements(1569) <= cp_elements(1568);
    -- CP-element group 1570 transition  bypass 
    -- predecessors 1568 
    -- successors 1571 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/ca
      -- 
    cp_elements(1570) <= cp_elements(1568);
    -- CP-element group 1571 join  transition  bypass 
    -- predecessors 1569 1570 
    -- successors 1578 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$exit
      -- 
    cp_element_group_1571: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1571"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1569) & cp_elements(1570);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1571), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1572 fork  transition  bypass 
    -- predecessors 1567 
    -- successors 1573 1575 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$entry
      -- 
    cp_elements(1572) <= cp_elements(1567);
    -- CP-element group 1573 transition  output  bypass 
    -- predecessors 1572 
    -- successors 1574 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/rr
      -- 
    cp_elements(1573) <= cp_elements(1572);
    rr_14853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1573), ack => type_cast_2508_inst_req_0); -- 
    -- CP-element group 1574 transition  input  bypass 
    -- predecessors 1573 
    -- successors 1577 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/ra
      -- 
    ra_14854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => cp_elements(1574)); -- 
    -- CP-element group 1575 transition  output  bypass 
    -- predecessors 1572 
    -- successors 1576 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/cr
      -- 
    cp_elements(1575) <= cp_elements(1572);
    cr_14858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1575), ack => type_cast_2508_inst_req_1); -- 
    -- CP-element group 1576 transition  input  bypass 
    -- predecessors 1575 
    -- successors 1577 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/ca
      -- 
    ca_14859_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => cp_elements(1576)); -- 
    -- CP-element group 1577 join  transition  bypass 
    -- predecessors 1574 1576 
    -- successors 1578 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$exit
      -- 
    cp_element_group_1577: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1577"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1574) & cp_elements(1576);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1577), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1578 join  transition  output  bypass 
    -- predecessors 1571 1577 
    -- successors 1583 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    cp_element_group_1578: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1578"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1571) & cp_elements(1577);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1578), clk => clk, reset => reset); --
    end block;
    phi_stmt_2503_req_14860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1578), ack => phi_stmt_2503_req_1); -- 
    -- CP-element group 1579 fork  transition  bypass 
    -- predecessors 1566 
    -- successors 1580 1581 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$entry
      -- 
    cp_elements(1579) <= cp_elements(1566);
    -- CP-element group 1580 transition  bypass 
    -- predecessors 1579 
    -- successors 1582 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/ra
      -- 
    cp_elements(1580) <= cp_elements(1579);
    -- CP-element group 1581 transition  bypass 
    -- predecessors 1579 
    -- successors 1582 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/ca
      -- 
    cp_elements(1581) <= cp_elements(1579);
    -- CP-element group 1582 join  transition  output  bypass 
    -- predecessors 1580 1581 
    -- successors 1583 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    cp_element_group_1582: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1582"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1580) & cp_elements(1581);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1582), clk => clk, reset => reset); --
    end block;
    phi_stmt_2509_req_14883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1582), ack => phi_stmt_2509_req_1); -- 
    -- CP-element group 1583 join  transition  bypass 
    -- predecessors 1578 1582 
    -- successors 1604 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xix_xpreheader_bbx_xnph7x_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1583: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1583"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1578) & cp_elements(1582);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1583), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1584 fork  transition  bypass 
    -- predecessors 666 
    -- successors 1585 1597 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1584) <= cp_elements(666);
    -- CP-element group 1585 fork  transition  bypass 
    -- predecessors 1584 
    -- successors 1586 1592 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- 
    cp_elements(1585) <= cp_elements(1584);
    -- CP-element group 1586 fork  transition  bypass 
    -- predecessors 1585 
    -- successors 1587 1589 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$entry
      -- 
    cp_elements(1586) <= cp_elements(1585);
    -- CP-element group 1587 transition  output  bypass 
    -- predecessors 1586 
    -- successors 1588 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/rr
      -- 
    cp_elements(1587) <= cp_elements(1586);
    rr_14902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1587), ack => type_cast_2506_inst_req_0); -- 
    -- CP-element group 1588 transition  input  bypass 
    -- predecessors 1587 
    -- successors 1591 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/ra
      -- 
    ra_14903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_0, ack => cp_elements(1588)); -- 
    -- CP-element group 1589 transition  output  bypass 
    -- predecessors 1586 
    -- successors 1590 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/cr
      -- 
    cp_elements(1589) <= cp_elements(1586);
    cr_14907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1589), ack => type_cast_2506_inst_req_1); -- 
    -- CP-element group 1590 transition  input  bypass 
    -- predecessors 1589 
    -- successors 1591 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/ca
      -- 
    ca_14908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_1, ack => cp_elements(1590)); -- 
    -- CP-element group 1591 join  transition  bypass 
    -- predecessors 1588 1590 
    -- successors 1596 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$exit
      -- 
    cp_element_group_1591: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1591"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1588) & cp_elements(1590);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1591), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1592 fork  transition  bypass 
    -- predecessors 1585 
    -- successors 1593 1594 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$entry
      -- 
    cp_elements(1592) <= cp_elements(1585);
    -- CP-element group 1593 transition  bypass 
    -- predecessors 1592 
    -- successors 1595 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/ra
      -- 
    cp_elements(1593) <= cp_elements(1592);
    -- CP-element group 1594 transition  bypass 
    -- predecessors 1592 
    -- successors 1595 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/ca
      -- 
    cp_elements(1594) <= cp_elements(1592);
    -- CP-element group 1595 join  transition  bypass 
    -- predecessors 1593 1594 
    -- successors 1596 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$exit
      -- 
    cp_element_group_1595: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1595"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1593) & cp_elements(1594);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1595), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1596 join  transition  output  bypass 
    -- predecessors 1591 1595 
    -- successors 1603 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    cp_element_group_1596: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1596"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1591) & cp_elements(1595);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1596), clk => clk, reset => reset); --
    end block;
    phi_stmt_2503_req_14925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1596), ack => phi_stmt_2503_req_0); -- 
    -- CP-element group 1597 fork  transition  bypass 
    -- predecessors 1584 
    -- successors 1598 1600 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$entry
      -- 
    cp_elements(1597) <= cp_elements(1584);
    -- CP-element group 1598 transition  output  bypass 
    -- predecessors 1597 
    -- successors 1599 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/rr
      -- 
    cp_elements(1598) <= cp_elements(1597);
    rr_14941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1598), ack => type_cast_2512_inst_req_0); -- 
    -- CP-element group 1599 transition  input  bypass 
    -- predecessors 1598 
    -- successors 1602 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/ra
      -- 
    ra_14942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_0, ack => cp_elements(1599)); -- 
    -- CP-element group 1600 transition  output  bypass 
    -- predecessors 1597 
    -- successors 1601 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/cr
      -- 
    cp_elements(1600) <= cp_elements(1597);
    cr_14946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1600), ack => type_cast_2512_inst_req_1); -- 
    -- CP-element group 1601 transition  input  bypass 
    -- predecessors 1600 
    -- successors 1602 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/ca
      -- 
    ca_14947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_1, ack => cp_elements(1601)); -- 
    -- CP-element group 1602 join  transition  output  bypass 
    -- predecessors 1599 1601 
    -- successors 1603 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    cp_element_group_1602: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1602"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1599) & cp_elements(1601);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1602), clk => clk, reset => reset); --
    end block;
    phi_stmt_2509_req_14948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1602), ack => phi_stmt_2509_req_0); -- 
    -- CP-element group 1603 join  transition  bypass 
    -- predecessors 1596 1602 
    -- successors 1604 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_bbx_xnph7x_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1603: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1603"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1596) & cp_elements(1602);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1603), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1604 merge  place  bypass 
    -- predecessors 1583 1603 
    -- successors 1605 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2502_PhiReqMerge
      -- 
    cp_elements(1604) <= OrReduce(cp_elements(1583) & cp_elements(1603));
    -- CP-element group 1605 fork  transition  bypass 
    -- predecessors 1604 
    -- successors 1606 1607 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2502_PhiAck/$entry
      -- 
    cp_elements(1605) <= cp_elements(1604);
    -- CP-element group 1606 transition  input  bypass 
    -- predecessors 1605 
    -- successors 1608 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2502_PhiAck/phi_stmt_2503_ack
      -- 
    phi_stmt_2503_ack_14953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2503_ack_0, ack => cp_elements(1606)); -- 
    -- CP-element group 1607 transition  input  bypass 
    -- predecessors 1605 
    -- successors 1608 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2502_PhiAck/phi_stmt_2509_ack
      -- 
    phi_stmt_2509_ack_14954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2509_ack_0, ack => cp_elements(1607)); -- 
    -- CP-element group 1608 join  transition  bypass 
    -- predecessors 1606 1607 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2502_PhiAck/$exit
      -- 
    cp_element_group_1608: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1608"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1606) & cp_elements(1607);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1608), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1609 fork  transition  bypass 
    -- predecessors 638 
    -- successors 1610 1622 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1609) <= cp_elements(638);
    -- CP-element group 1610 fork  transition  bypass 
    -- predecessors 1609 
    -- successors 1611 1617 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/$entry
      -- 
    cp_elements(1610) <= cp_elements(1609);
    -- CP-element group 1611 fork  transition  bypass 
    -- predecessors 1610 
    -- successors 1612 1614 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/$entry
      -- 
    cp_elements(1611) <= cp_elements(1610);
    -- CP-element group 1612 transition  output  bypass 
    -- predecessors 1611 
    -- successors 1613 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/rr
      -- 
    cp_elements(1612) <= cp_elements(1611);
    rr_14985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1612), ack => type_cast_2540_inst_req_0); -- 
    -- CP-element group 1613 transition  input  bypass 
    -- predecessors 1612 
    -- successors 1616 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/ra
      -- 
    ra_14986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2540_inst_ack_0, ack => cp_elements(1613)); -- 
    -- CP-element group 1614 transition  output  bypass 
    -- predecessors 1611 
    -- successors 1615 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/cr
      -- 
    cp_elements(1614) <= cp_elements(1611);
    cr_14990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1614), ack => type_cast_2540_inst_req_1); -- 
    -- CP-element group 1615 transition  input  bypass 
    -- predecessors 1614 
    -- successors 1616 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/ca
      -- 
    ca_14991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2540_inst_ack_1, ack => cp_elements(1615)); -- 
    -- CP-element group 1616 join  transition  bypass 
    -- predecessors 1613 1615 
    -- successors 1621 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/$exit
      -- 
    cp_element_group_1616: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1616"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1613) & cp_elements(1615);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1616), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1617 fork  transition  bypass 
    -- predecessors 1610 
    -- successors 1618 1619 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/$entry
      -- 
    cp_elements(1617) <= cp_elements(1610);
    -- CP-element group 1618 transition  bypass 
    -- predecessors 1617 
    -- successors 1620 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/ra
      -- 
    cp_elements(1618) <= cp_elements(1617);
    -- CP-element group 1619 transition  bypass 
    -- predecessors 1617 
    -- successors 1620 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/ca
      -- 
    cp_elements(1619) <= cp_elements(1617);
    -- CP-element group 1620 join  transition  bypass 
    -- predecessors 1618 1619 
    -- successors 1621 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/$exit
      -- 
    cp_element_group_1620: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1620"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1618) & cp_elements(1619);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1620), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1621 join  transition  output  bypass 
    -- predecessors 1616 1620 
    -- successors 1628 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_req
      -- 
    cp_element_group_1621: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1621"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1616) & cp_elements(1620);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1621), clk => clk, reset => reset); --
    end block;
    phi_stmt_2537_req_15008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1621), ack => phi_stmt_2537_req_0); -- 
    -- CP-element group 1622 fork  transition  bypass 
    -- predecessors 1609 
    -- successors 1623 1625 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$entry
      -- 
    cp_elements(1622) <= cp_elements(1609);
    -- CP-element group 1623 transition  output  bypass 
    -- predecessors 1622 
    -- successors 1624 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/rr
      -- 
    cp_elements(1623) <= cp_elements(1622);
    rr_15024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1623), ack => type_cast_2546_inst_req_0); -- 
    -- CP-element group 1624 transition  input  bypass 
    -- predecessors 1623 
    -- successors 1627 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/ra
      -- 
    ra_15025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_0, ack => cp_elements(1624)); -- 
    -- CP-element group 1625 transition  output  bypass 
    -- predecessors 1622 
    -- successors 1626 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/cr
      -- 
    cp_elements(1625) <= cp_elements(1622);
    cr_15029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1625), ack => type_cast_2546_inst_req_1); -- 
    -- CP-element group 1626 transition  input  bypass 
    -- predecessors 1625 
    -- successors 1627 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/ca
      -- 
    ca_15030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_1, ack => cp_elements(1626)); -- 
    -- CP-element group 1627 join  transition  output  bypass 
    -- predecessors 1624 1626 
    -- successors 1628 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_req
      -- 
    cp_element_group_1627: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1627"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1624) & cp_elements(1626);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1627), clk => clk, reset => reset); --
    end block;
    phi_stmt_2543_req_15031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1627), ack => phi_stmt_2543_req_0); -- 
    -- CP-element group 1628 join  transition  bypass 
    -- predecessors 1621 1627 
    -- successors 1647 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_bbx_xnphx_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1628: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1628"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1621) & cp_elements(1627);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1628), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1629 fork  transition  bypass 
    -- predecessors 31 
    -- successors 1630 1642 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1629) <= cp_elements(31);
    -- CP-element group 1630 fork  transition  bypass 
    -- predecessors 1629 
    -- successors 1631 1635 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/$entry
      -- 
    cp_elements(1630) <= cp_elements(1629);
    -- CP-element group 1631 fork  transition  bypass 
    -- predecessors 1630 
    -- successors 1632 1633 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/$entry
      -- 
    cp_elements(1631) <= cp_elements(1630);
    -- CP-element group 1632 transition  bypass 
    -- predecessors 1631 
    -- successors 1634 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Sample/ra
      -- 
    cp_elements(1632) <= cp_elements(1631);
    -- CP-element group 1633 transition  bypass 
    -- predecessors 1631 
    -- successors 1634 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/Update/ca
      -- 
    cp_elements(1633) <= cp_elements(1631);
    -- CP-element group 1634 join  transition  bypass 
    -- predecessors 1632 1633 
    -- successors 1641 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2540/SplitProtocol/$exit
      -- 
    cp_element_group_1634: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1634"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1632) & cp_elements(1633);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1634), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1635 fork  transition  bypass 
    -- predecessors 1630 
    -- successors 1636 1638 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/$entry
      -- 
    cp_elements(1635) <= cp_elements(1630);
    -- CP-element group 1636 transition  output  bypass 
    -- predecessors 1635 
    -- successors 1637 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/rr
      -- 
    cp_elements(1636) <= cp_elements(1635);
    rr_15066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1636), ack => type_cast_2542_inst_req_0); -- 
    -- CP-element group 1637 transition  input  bypass 
    -- predecessors 1636 
    -- successors 1640 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Sample/ra
      -- 
    ra_15067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2542_inst_ack_0, ack => cp_elements(1637)); -- 
    -- CP-element group 1638 transition  output  bypass 
    -- predecessors 1635 
    -- successors 1639 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/cr
      -- 
    cp_elements(1638) <= cp_elements(1635);
    cr_15071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1638), ack => type_cast_2542_inst_req_1); -- 
    -- CP-element group 1639 transition  input  bypass 
    -- predecessors 1638 
    -- successors 1640 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/Update/ca
      -- 
    ca_15072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2542_inst_ack_1, ack => cp_elements(1639)); -- 
    -- CP-element group 1640 join  transition  bypass 
    -- predecessors 1637 1639 
    -- successors 1641 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/type_cast_2542/SplitProtocol/$exit
      -- 
    cp_element_group_1640: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1640"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1637) & cp_elements(1639);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1640), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1641 join  transition  output  bypass 
    -- predecessors 1634 1640 
    -- successors 1646 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2537/phi_stmt_2537_req
      -- 
    cp_element_group_1641: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1641"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1634) & cp_elements(1640);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1641), clk => clk, reset => reset); --
    end block;
    phi_stmt_2537_req_15073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1641), ack => phi_stmt_2537_req_1); -- 
    -- CP-element group 1642 fork  transition  bypass 
    -- predecessors 1629 
    -- successors 1643 1644 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$entry
      -- 
    cp_elements(1642) <= cp_elements(1629);
    -- CP-element group 1643 transition  bypass 
    -- predecessors 1642 
    -- successors 1645 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/ra
      -- 
    cp_elements(1643) <= cp_elements(1642);
    -- CP-element group 1644 transition  bypass 
    -- predecessors 1642 
    -- successors 1645 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/ca
      -- 
    cp_elements(1644) <= cp_elements(1642);
    -- CP-element group 1645 join  transition  output  bypass 
    -- predecessors 1643 1644 
    -- successors 1646 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/phi_stmt_2543/phi_stmt_2543_req
      -- 
    cp_element_group_1645: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1645"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1643) & cp_elements(1644);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1645), clk => clk, reset => reset); --
    end block;
    phi_stmt_2543_req_15096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1645), ack => phi_stmt_2543_req_1); -- 
    -- CP-element group 1646 join  transition  bypass 
    -- predecessors 1641 1645 
    -- successors 1647 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xix_xpreheader_bbx_xnphx_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1646: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1646"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1641) & cp_elements(1645);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1646), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1647 merge  place  bypass 
    -- predecessors 1628 1646 
    -- successors 1648 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2536_PhiReqMerge
      -- 
    cp_elements(1647) <= OrReduce(cp_elements(1628) & cp_elements(1646));
    -- CP-element group 1648 fork  transition  bypass 
    -- predecessors 1647 
    -- successors 1649 1650 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2536_PhiAck/$entry
      -- 
    cp_elements(1648) <= cp_elements(1647);
    -- CP-element group 1649 transition  input  bypass 
    -- predecessors 1648 
    -- successors 1651 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2536_PhiAck/phi_stmt_2537_ack
      -- 
    phi_stmt_2537_ack_15101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2537_ack_0, ack => cp_elements(1649)); -- 
    -- CP-element group 1650 transition  input  bypass 
    -- predecessors 1648 
    -- successors 1651 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2536_PhiAck/phi_stmt_2543_ack
      -- 
    phi_stmt_2543_ack_15102_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2543_ack_0, ack => cp_elements(1650)); -- 
    -- CP-element group 1651 join  transition  bypass 
    -- predecessors 1649 1650 
    -- successors 32 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2536_PhiAck/$exit
      -- 
    cp_element_group_1651: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1651"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1649) & cp_elements(1650);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1651), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1652 fork  transition  bypass 
    -- predecessors 640 
    -- successors 1653 1659 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/$entry
      -- 
    cp_elements(1652) <= cp_elements(640);
    -- CP-element group 1653 fork  transition  bypass 
    -- predecessors 1652 
    -- successors 1654 1656 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/$entry
      -- 
    cp_elements(1653) <= cp_elements(1652);
    -- CP-element group 1654 transition  output  bypass 
    -- predecessors 1653 
    -- successors 1655 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Sample/rr
      -- 
    cp_elements(1654) <= cp_elements(1653);
    rr_15125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1654), ack => type_cast_2578_inst_req_0); -- 
    -- CP-element group 1655 transition  input  bypass 
    -- predecessors 1654 
    -- successors 1658 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Sample/ra
      -- 
    ra_15126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2578_inst_ack_0, ack => cp_elements(1655)); -- 
    -- CP-element group 1656 transition  output  bypass 
    -- predecessors 1653 
    -- successors 1657 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Update/cr
      -- 
    cp_elements(1656) <= cp_elements(1653);
    cr_15130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1656), ack => type_cast_2578_inst_req_1); -- 
    -- CP-element group 1657 transition  input  bypass 
    -- predecessors 1656 
    -- successors 1658 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/Update/ca
      -- 
    ca_15131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2578_inst_ack_1, ack => cp_elements(1657)); -- 
    -- CP-element group 1658 join  transition  output  bypass 
    -- predecessors 1655 1657 
    -- successors 1665 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_sources/type_cast_2578/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2575/phi_stmt_2575_req
      -- 
    cp_element_group_1658: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1658"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1655) & cp_elements(1657);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1658), clk => clk, reset => reset); --
    end block;
    phi_stmt_2575_req_15132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1658), ack => phi_stmt_2575_req_0); -- 
    -- CP-element group 1659 fork  transition  bypass 
    -- predecessors 1652 
    -- successors 1660 1662 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/$entry
      -- 
    cp_elements(1659) <= cp_elements(1652);
    -- CP-element group 1660 transition  output  bypass 
    -- predecessors 1659 
    -- successors 1661 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Sample/rr
      -- 
    cp_elements(1660) <= cp_elements(1659);
    rr_15148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1660), ack => type_cast_2582_inst_req_0); -- 
    -- CP-element group 1661 transition  input  bypass 
    -- predecessors 1660 
    -- successors 1664 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Sample/ra
      -- 
    ra_15149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_0, ack => cp_elements(1661)); -- 
    -- CP-element group 1662 transition  output  bypass 
    -- predecessors 1659 
    -- successors 1663 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Update/cr
      -- 
    cp_elements(1662) <= cp_elements(1659);
    cr_15153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1662), ack => type_cast_2582_inst_req_1); -- 
    -- CP-element group 1663 transition  input  bypass 
    -- predecessors 1662 
    -- successors 1664 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/Update/ca
      -- 
    ca_15154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_1, ack => cp_elements(1663)); -- 
    -- CP-element group 1664 join  transition  output  bypass 
    -- predecessors 1661 1663 
    -- successors 1665 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_sources/type_cast_2582/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2579/phi_stmt_2579_req
      -- 
    cp_element_group_1664: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1664"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1661) & cp_elements(1663);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1664), clk => clk, reset => reset); --
    end block;
    phi_stmt_2579_req_15155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1664), ack => phi_stmt_2579_req_0); -- 
    -- CP-element group 1665 join  transition  bypass 
    -- predecessors 1658 1664 
    -- successors 1666 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xi_xx_x_crit_edgex_xix_xix_xix_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_1665: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1665"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1658) & cp_elements(1664);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1665), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1666 place  bypass 
    -- predecessors 1665 
    -- successors 1667 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2574_PhiReqMerge
      -- 
    cp_elements(1666) <= cp_elements(1665);
    -- CP-element group 1667 fork  transition  bypass 
    -- predecessors 1666 
    -- successors 1668 1669 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2574_PhiAck/$entry
      -- 
    cp_elements(1667) <= cp_elements(1666);
    -- CP-element group 1668 transition  input  bypass 
    -- predecessors 1667 
    -- successors 1670 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2574_PhiAck/phi_stmt_2575_ack
      -- 
    phi_stmt_2575_ack_15160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2575_ack_0, ack => cp_elements(1668)); -- 
    -- CP-element group 1669 transition  input  bypass 
    -- predecessors 1667 
    -- successors 1670 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2574_PhiAck/phi_stmt_2579_ack
      -- 
    phi_stmt_2579_ack_15161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2579_ack_0, ack => cp_elements(1669)); -- 
    -- CP-element group 1670 join  transition  bypass 
    -- predecessors 1668 1669 
    -- successors 34 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2574_PhiAck/$exit
      -- 
    cp_element_group_1670: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1670"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1668) & cp_elements(1669);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1670), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1671 fork  transition  bypass 
    -- predecessors 618 
    -- successors 1672 1684 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1671) <= cp_elements(618);
    -- CP-element group 1672 fork  transition  bypass 
    -- predecessors 1671 
    -- successors 1673 1679 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/$entry
      -- 
    cp_elements(1672) <= cp_elements(1671);
    -- CP-element group 1673 fork  transition  bypass 
    -- predecessors 1672 
    -- successors 1674 1676 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/$entry
      -- 
    cp_elements(1673) <= cp_elements(1672);
    -- CP-element group 1674 transition  output  bypass 
    -- predecessors 1673 
    -- successors 1675 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/rr
      -- 
    cp_elements(1674) <= cp_elements(1673);
    rr_15180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1674), ack => type_cast_2589_inst_req_0); -- 
    -- CP-element group 1675 transition  input  bypass 
    -- predecessors 1674 
    -- successors 1678 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/ra
      -- 
    ra_15181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_0, ack => cp_elements(1675)); -- 
    -- CP-element group 1676 transition  output  bypass 
    -- predecessors 1673 
    -- successors 1677 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/cr
      -- 
    cp_elements(1676) <= cp_elements(1673);
    cr_15185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1676), ack => type_cast_2589_inst_req_1); -- 
    -- CP-element group 1677 transition  input  bypass 
    -- predecessors 1676 
    -- successors 1678 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/ca
      -- 
    ca_15186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_1, ack => cp_elements(1677)); -- 
    -- CP-element group 1678 join  transition  bypass 
    -- predecessors 1675 1677 
    -- successors 1683 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/$exit
      -- 
    cp_element_group_1678: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1678"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1675) & cp_elements(1677);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1678), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1679 fork  transition  bypass 
    -- predecessors 1672 
    -- successors 1680 1681 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/$entry
      -- 
    cp_elements(1679) <= cp_elements(1672);
    -- CP-element group 1680 transition  bypass 
    -- predecessors 1679 
    -- successors 1682 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/ra
      -- 
    cp_elements(1680) <= cp_elements(1679);
    -- CP-element group 1681 transition  bypass 
    -- predecessors 1679 
    -- successors 1682 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/ca
      -- 
    cp_elements(1681) <= cp_elements(1679);
    -- CP-element group 1682 join  transition  bypass 
    -- predecessors 1680 1681 
    -- successors 1683 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/$exit
      -- 
    cp_element_group_1682: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1682"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1680) & cp_elements(1681);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1682), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1683 join  transition  output  bypass 
    -- predecessors 1678 1682 
    -- successors 1688 
    -- members (3) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_req
      -- 
    cp_element_group_1683: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1683"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1678) & cp_elements(1682);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1683), clk => clk, reset => reset); --
    end block;
    phi_stmt_2586_req_15203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1683), ack => phi_stmt_2586_req_0); -- 
    -- CP-element group 1684 fork  transition  bypass 
    -- predecessors 1671 
    -- successors 1685 1686 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/$entry
      -- 
    cp_elements(1684) <= cp_elements(1671);
    -- CP-element group 1685 transition  bypass 
    -- predecessors 1684 
    -- successors 1687 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/ra
      -- 
    cp_elements(1685) <= cp_elements(1684);
    -- CP-element group 1686 transition  bypass 
    -- predecessors 1684 
    -- successors 1687 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/ca
      -- 
    cp_elements(1686) <= cp_elements(1684);
    -- CP-element group 1687 join  transition  output  bypass 
    -- predecessors 1685 1686 
    -- successors 1688 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_req
      -- 
    cp_element_group_1687: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1687"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1685) & cp_elements(1686);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1687), clk => clk, reset => reset); --
    end block;
    phi_stmt_2592_req_15226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1687), ack => phi_stmt_2592_req_0); -- 
    -- CP-element group 1688 join  transition  bypass 
    -- predecessors 1683 1687 
    -- successors 1709 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xix_xi_xx_x_crit_edgex_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1688: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1688"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1683) & cp_elements(1687);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1688), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1689 fork  transition  bypass 
    -- predecessors 34 
    -- successors 1690 1702 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1689) <= cp_elements(34);
    -- CP-element group 1690 fork  transition  bypass 
    -- predecessors 1689 
    -- successors 1691 1695 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/$entry
      -- 
    cp_elements(1690) <= cp_elements(1689);
    -- CP-element group 1691 fork  transition  bypass 
    -- predecessors 1690 
    -- successors 1692 1693 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/$entry
      -- 
    cp_elements(1691) <= cp_elements(1690);
    -- CP-element group 1692 transition  bypass 
    -- predecessors 1691 
    -- successors 1694 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Sample/ra
      -- 
    cp_elements(1692) <= cp_elements(1691);
    -- CP-element group 1693 transition  bypass 
    -- predecessors 1691 
    -- successors 1694 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/Update/ca
      -- 
    cp_elements(1693) <= cp_elements(1691);
    -- CP-element group 1694 join  transition  bypass 
    -- predecessors 1692 1693 
    -- successors 1701 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2589/SplitProtocol/$exit
      -- 
    cp_element_group_1694: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1694"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1692) & cp_elements(1693);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1694), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1695 fork  transition  bypass 
    -- predecessors 1690 
    -- successors 1696 1698 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/$entry
      -- 
    cp_elements(1695) <= cp_elements(1690);
    -- CP-element group 1696 transition  output  bypass 
    -- predecessors 1695 
    -- successors 1697 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/rr
      -- 
    cp_elements(1696) <= cp_elements(1695);
    rr_15261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1696), ack => type_cast_2591_inst_req_0); -- 
    -- CP-element group 1697 transition  input  bypass 
    -- predecessors 1696 
    -- successors 1700 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Sample/ra
      -- 
    ra_15262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_0, ack => cp_elements(1697)); -- 
    -- CP-element group 1698 transition  output  bypass 
    -- predecessors 1695 
    -- successors 1699 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/cr
      -- 
    cp_elements(1698) <= cp_elements(1695);
    cr_15266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1698), ack => type_cast_2591_inst_req_1); -- 
    -- CP-element group 1699 transition  input  bypass 
    -- predecessors 1698 
    -- successors 1700 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/Update/ca
      -- 
    ca_15267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_1, ack => cp_elements(1699)); -- 
    -- CP-element group 1700 join  transition  bypass 
    -- predecessors 1697 1699 
    -- successors 1701 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/type_cast_2591/SplitProtocol/$exit
      -- 
    cp_element_group_1700: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1700"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1697) & cp_elements(1699);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1700), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1701 join  transition  output  bypass 
    -- predecessors 1694 1700 
    -- successors 1708 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2586/phi_stmt_2586_req
      -- 
    cp_element_group_1701: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1701"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1694) & cp_elements(1700);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1701), clk => clk, reset => reset); --
    end block;
    phi_stmt_2586_req_15268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1701), ack => phi_stmt_2586_req_1); -- 
    -- CP-element group 1702 fork  transition  bypass 
    -- predecessors 1689 
    -- successors 1703 1705 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/$entry
      -- 
    cp_elements(1702) <= cp_elements(1689);
    -- CP-element group 1703 transition  output  bypass 
    -- predecessors 1702 
    -- successors 1704 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/rr
      -- 
    cp_elements(1703) <= cp_elements(1702);
    rr_15284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1703), ack => type_cast_2598_inst_req_0); -- 
    -- CP-element group 1704 transition  input  bypass 
    -- predecessors 1703 
    -- successors 1707 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Sample/ra
      -- 
    ra_15285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_0, ack => cp_elements(1704)); -- 
    -- CP-element group 1705 transition  output  bypass 
    -- predecessors 1702 
    -- successors 1706 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/cr
      -- 
    cp_elements(1705) <= cp_elements(1702);
    cr_15289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1705), ack => type_cast_2598_inst_req_1); -- 
    -- CP-element group 1706 transition  input  bypass 
    -- predecessors 1705 
    -- successors 1707 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/Update/ca
      -- 
    ca_15290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_1, ack => cp_elements(1706)); -- 
    -- CP-element group 1707 join  transition  output  bypass 
    -- predecessors 1704 1706 
    -- successors 1708 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_sources/type_cast_2598/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/phi_stmt_2592/phi_stmt_2592_req
      -- 
    cp_element_group_1707: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1707"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1704) & cp_elements(1706);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1707), clk => clk, reset => reset); --
    end block;
    phi_stmt_2592_req_15291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1707), ack => phi_stmt_2592_req_1); -- 
    -- CP-element group 1708 join  transition  bypass 
    -- predecessors 1701 1707 
    -- successors 1709 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xix_xloopexit_xx_x_crit_edgex_xix_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1708: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1708"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1701) & cp_elements(1707);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1708), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1709 merge  place  bypass 
    -- predecessors 1688 1708 
    -- successors 1710 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2585_PhiReqMerge
      -- 
    cp_elements(1709) <= OrReduce(cp_elements(1688) & cp_elements(1708));
    -- CP-element group 1710 fork  transition  bypass 
    -- predecessors 1709 
    -- successors 1711 1712 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2585_PhiAck/$entry
      -- 
    cp_elements(1710) <= cp_elements(1709);
    -- CP-element group 1711 transition  input  bypass 
    -- predecessors 1710 
    -- successors 1713 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2585_PhiAck/phi_stmt_2586_ack
      -- 
    phi_stmt_2586_ack_15296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2586_ack_0, ack => cp_elements(1711)); -- 
    -- CP-element group 1712 transition  input  bypass 
    -- predecessors 1710 
    -- successors 1713 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2585_PhiAck/phi_stmt_2592_ack
      -- 
    phi_stmt_2592_ack_15297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2592_ack_0, ack => cp_elements(1712)); -- 
    -- CP-element group 1713 join  transition  bypass 
    -- predecessors 1711 1712 
    -- successors 35 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2585_PhiAck/$exit
      -- 
    cp_element_group_1713: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1713"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1711) & cp_elements(1712);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1713), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1714 transition  output  bypass 
    -- predecessors 664 
    -- successors 1715 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Sample/rr
      -- 
    cp_elements(1714) <= cp_elements(664);
    rr_15320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1714), ack => type_cast_2625_inst_req_0); -- 
    -- CP-element group 1715 transition  input  bypass 
    -- predecessors 1714 
    -- successors 1718 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Sample/ra
      -- 
    ra_15321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2625_inst_ack_0, ack => cp_elements(1715)); -- 
    -- CP-element group 1716 transition  output  bypass 
    -- predecessors 664 
    -- successors 1717 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Update/cr
      -- 
    cp_elements(1716) <= cp_elements(664);
    cr_15325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1716), ack => type_cast_2625_inst_req_1); -- 
    -- CP-element group 1717 transition  input  bypass 
    -- predecessors 1716 
    -- successors 1718 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/Update/ca
      -- 
    ca_15326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2625_inst_ack_1, ack => cp_elements(1717)); -- 
    -- CP-element group 1718 join  transition  place  output  bypass 
    -- predecessors 1715 1717 
    -- successors 1719 
    -- members (8) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_sources/type_cast_2625/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xi_xx_xloopexitx_xix_xix_xix_xloopexit_PhiReq/phi_stmt_2622/phi_stmt_2622_req
      -- 	branch_block_stmt_1659/merge_stmt_2621_PhiReqMerge
      -- 	branch_block_stmt_1659/merge_stmt_2621_PhiAck/$entry
      -- 
    cp_element_group_1718: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1718"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1715) & cp_elements(1717);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1718), clk => clk, reset => reset); --
    end block;
    phi_stmt_2622_req_15327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1718), ack => phi_stmt_2622_req_0); -- 
    -- CP-element group 1719 transition  input  bypass 
    -- predecessors 1718 
    -- successors 37 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2621_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2621_PhiAck/phi_stmt_2622_ack
      -- 
    phi_stmt_2622_ack_15332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2622_ack_0, ack => cp_elements(1719)); -- 
    -- CP-element group 1720 transition  bypass 
    -- predecessors 597 
    -- successors 1722 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/ra
      -- 
    cp_elements(1720) <= cp_elements(597);
    -- CP-element group 1721 transition  bypass 
    -- predecessors 597 
    -- successors 1722 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/ca
      -- 
    cp_elements(1721) <= cp_elements(597);
    -- CP-element group 1722 join  transition  output  bypass 
    -- predecessors 1720 1721 
    -- successors 1728 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_27_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_req
      -- 
    cp_element_group_1722: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1722"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1720) & cp_elements(1721);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1722), clk => clk, reset => reset); --
    end block;
    phi_stmt_2629_req_15358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1722), ack => phi_stmt_2629_req_0); -- 
    -- CP-element group 1723 transition  output  bypass 
    -- predecessors 37 
    -- successors 1724 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/rr
      -- 
    cp_elements(1723) <= cp_elements(37);
    rr_15377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1723), ack => type_cast_2635_inst_req_0); -- 
    -- CP-element group 1724 transition  input  bypass 
    -- predecessors 1723 
    -- successors 1727 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Sample/ra
      -- 
    ra_15378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2635_inst_ack_0, ack => cp_elements(1724)); -- 
    -- CP-element group 1725 transition  output  bypass 
    -- predecessors 37 
    -- successors 1726 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/cr
      -- 
    cp_elements(1725) <= cp_elements(37);
    cr_15382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1725), ack => type_cast_2635_inst_req_1); -- 
    -- CP-element group 1726 transition  input  bypass 
    -- predecessors 1725 
    -- successors 1727 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/Update/ca
      -- 
    ca_15383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2635_inst_ack_1, ack => cp_elements(1726)); -- 
    -- CP-element group 1727 join  transition  output  bypass 
    -- predecessors 1724 1726 
    -- successors 1728 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_sources/type_cast_2635/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xix_xloopexit_xx_xloopexitx_xix_xix_xi_PhiReq/phi_stmt_2629/phi_stmt_2629_req
      -- 
    cp_element_group_1727: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1727"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1724) & cp_elements(1726);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1727), clk => clk, reset => reset); --
    end block;
    phi_stmt_2629_req_15384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1727), ack => phi_stmt_2629_req_1); -- 
    -- CP-element group 1728 merge  place  bypass 
    -- predecessors 1722 1727 
    -- successors 1729 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2628_PhiReqMerge
      -- 
    cp_elements(1728) <= OrReduce(cp_elements(1722) & cp_elements(1727));
    -- CP-element group 1729 transition  bypass 
    -- predecessors 1728 
    -- successors 1730 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2628_PhiAck/$entry
      -- 
    cp_elements(1729) <= cp_elements(1728);
    -- CP-element group 1730 fork  transition  place  input  bypass 
    -- predecessors 1729 
    -- successors 1742 1748 
    -- members (7) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi
      -- 	branch_block_stmt_1659/merge_stmt_2628__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2628_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2628_PhiAck/phi_stmt_2629_ack
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/$entry
      -- 
    phi_stmt_2629_ack_15389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2629_ack_0, ack => cp_elements(1730)); -- 
    -- CP-element group 1731 fork  transition  bypass 
    -- predecessors 599 
    -- successors 1732 1733 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/$entry
      -- 
    cp_elements(1731) <= cp_elements(599);
    -- CP-element group 1732 transition  bypass 
    -- predecessors 1731 
    -- successors 1734 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/ra
      -- 
    cp_elements(1732) <= cp_elements(1731);
    -- CP-element group 1733 transition  bypass 
    -- predecessors 1731 
    -- successors 1734 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/ca
      -- 
    cp_elements(1733) <= cp_elements(1731);
    -- CP-element group 1734 join  transition  bypass 
    -- predecessors 1732 1733 
    -- successors 1741 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/$exit
      -- 
    cp_element_group_1734: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1734"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1732) & cp_elements(1733);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1734), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1735 fork  transition  bypass 
    -- predecessors 599 
    -- successors 1736 1738 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/$entry
      -- 
    cp_elements(1735) <= cp_elements(599);
    -- CP-element group 1736 transition  output  bypass 
    -- predecessors 1735 
    -- successors 1737 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/rr
      -- 
    cp_elements(1736) <= cp_elements(1735);
    rr_15424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1736), ack => type_cast_2644_inst_req_0); -- 
    -- CP-element group 1737 transition  input  bypass 
    -- predecessors 1736 
    -- successors 1740 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/ra
      -- 
    ra_15425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2644_inst_ack_0, ack => cp_elements(1737)); -- 
    -- CP-element group 1738 transition  output  bypass 
    -- predecessors 1735 
    -- successors 1739 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/cr
      -- 
    cp_elements(1738) <= cp_elements(1735);
    cr_15429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1738), ack => type_cast_2644_inst_req_1); -- 
    -- CP-element group 1739 transition  input  bypass 
    -- predecessors 1738 
    -- successors 1740 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/ca
      -- 
    ca_15430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2644_inst_ack_1, ack => cp_elements(1739)); -- 
    -- CP-element group 1740 join  transition  bypass 
    -- predecessors 1737 1739 
    -- successors 1741 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/$exit
      -- 
    cp_element_group_1740: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1740"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1737) & cp_elements(1739);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1740), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1741 join  transition  output  bypass 
    -- predecessors 1734 1740 
    -- successors 1753 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/$exit
      -- 	branch_block_stmt_1659/bb_27_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_req
      -- 
    cp_element_group_1741: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1741"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1734) & cp_elements(1740);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1741), clk => clk, reset => reset); --
    end block;
    phi_stmt_2639_req_15431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1741), ack => phi_stmt_2639_req_1); -- 
    -- CP-element group 1742 fork  transition  bypass 
    -- predecessors 1730 
    -- successors 1743 1745 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/$entry
      -- 
    cp_elements(1742) <= cp_elements(1730);
    -- CP-element group 1743 transition  output  bypass 
    -- predecessors 1742 
    -- successors 1744 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/rr
      -- 
    cp_elements(1743) <= cp_elements(1742);
    rr_15450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1743), ack => type_cast_2642_inst_req_0); -- 
    -- CP-element group 1744 transition  input  bypass 
    -- predecessors 1743 
    -- successors 1747 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Sample/ra
      -- 
    ra_15451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2642_inst_ack_0, ack => cp_elements(1744)); -- 
    -- CP-element group 1745 transition  output  bypass 
    -- predecessors 1742 
    -- successors 1746 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/cr
      -- 
    cp_elements(1745) <= cp_elements(1742);
    cr_15455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1745), ack => type_cast_2642_inst_req_1); -- 
    -- CP-element group 1746 transition  input  bypass 
    -- predecessors 1745 
    -- successors 1747 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/Update/ca
      -- 
    ca_15456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2642_inst_ack_1, ack => cp_elements(1746)); -- 
    -- CP-element group 1747 join  transition  bypass 
    -- predecessors 1744 1746 
    -- successors 1752 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2642/SplitProtocol/$exit
      -- 
    cp_element_group_1747: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1747"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1744) & cp_elements(1746);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1747), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1748 fork  transition  bypass 
    -- predecessors 1730 
    -- successors 1749 1750 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/$entry
      -- 
    cp_elements(1748) <= cp_elements(1730);
    -- CP-element group 1749 transition  bypass 
    -- predecessors 1748 
    -- successors 1751 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Sample/ra
      -- 
    cp_elements(1749) <= cp_elements(1748);
    -- CP-element group 1750 transition  bypass 
    -- predecessors 1748 
    -- successors 1751 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/Update/ca
      -- 
    cp_elements(1750) <= cp_elements(1748);
    -- CP-element group 1751 join  transition  bypass 
    -- predecessors 1749 1750 
    -- successors 1752 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/type_cast_2644/SplitProtocol/$exit
      -- 
    cp_element_group_1751: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1751"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1749) & cp_elements(1750);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1751), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1752 join  transition  output  bypass 
    -- predecessors 1747 1751 
    -- successors 1753 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_sources/$exit
      -- 	branch_block_stmt_1659/xx_xloopexitx_xix_xix_xi_udiv32x_xexitx_xpreheaderx_xix_xi_PhiReq/phi_stmt_2639/phi_stmt_2639_req
      -- 
    cp_element_group_1752: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1752"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1747) & cp_elements(1751);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1752), clk => clk, reset => reset); --
    end block;
    phi_stmt_2639_req_15473_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1752), ack => phi_stmt_2639_req_0); -- 
    -- CP-element group 1753 merge  place  bypass 
    -- predecessors 1741 1752 
    -- successors 1754 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2638_PhiReqMerge
      -- 
    cp_elements(1753) <= OrReduce(cp_elements(1741) & cp_elements(1752));
    -- CP-element group 1754 transition  bypass 
    -- predecessors 1753 
    -- successors 1755 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2638_PhiAck/$entry
      -- 
    cp_elements(1754) <= cp_elements(1753);
    -- CP-element group 1755 transition  place  input  bypass 
    -- predecessors 1754 
    -- successors 667 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2651_to_assign_stmt_2670__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2638__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2638_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2638_PhiAck/phi_stmt_2639_ack
      -- 
    phi_stmt_2639_ack_15478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2639_ack_0, ack => cp_elements(1755)); -- 
    -- CP-element group 1756 fork  transition  bypass 
    -- predecessors 723 
    -- successors 1757 1763 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1756) <= cp_elements(723);
    -- CP-element group 1757 fork  transition  bypass 
    -- predecessors 1756 
    -- successors 1758 1760 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/$entry
      -- 
    cp_elements(1757) <= cp_elements(1756);
    -- CP-element group 1758 transition  output  bypass 
    -- predecessors 1757 
    -- successors 1759 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/rr
      -- 
    cp_elements(1758) <= cp_elements(1757);
    rr_15509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1758), ack => type_cast_2683_inst_req_0); -- 
    -- CP-element group 1759 transition  input  bypass 
    -- predecessors 1758 
    -- successors 1762 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/ra
      -- 
    ra_15510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2683_inst_ack_0, ack => cp_elements(1759)); -- 
    -- CP-element group 1760 transition  output  bypass 
    -- predecessors 1757 
    -- successors 1761 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/cr
      -- 
    cp_elements(1760) <= cp_elements(1757);
    cr_15514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1760), ack => type_cast_2683_inst_req_1); -- 
    -- CP-element group 1761 transition  input  bypass 
    -- predecessors 1760 
    -- successors 1762 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/ca
      -- 
    ca_15515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2683_inst_ack_1, ack => cp_elements(1761)); -- 
    -- CP-element group 1762 join  transition  output  bypass 
    -- predecessors 1759 1761 
    -- successors 1775 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_req
      -- 
    cp_element_group_1762: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1762"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1759) & cp_elements(1761);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1762), clk => clk, reset => reset); --
    end block;
    phi_stmt_2680_req_15516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1762), ack => phi_stmt_2680_req_0); -- 
    -- CP-element group 1763 fork  transition  bypass 
    -- predecessors 1756 
    -- successors 1764 1770 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/$entry
      -- 
    cp_elements(1763) <= cp_elements(1756);
    -- CP-element group 1764 fork  transition  bypass 
    -- predecessors 1763 
    -- successors 1765 1767 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/$entry
      -- 
    cp_elements(1764) <= cp_elements(1763);
    -- CP-element group 1765 transition  output  bypass 
    -- predecessors 1764 
    -- successors 1766 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/rr
      -- 
    cp_elements(1765) <= cp_elements(1764);
    rr_15532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1765), ack => type_cast_2690_inst_req_0); -- 
    -- CP-element group 1766 transition  input  bypass 
    -- predecessors 1765 
    -- successors 1769 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/ra
      -- 
    ra_15533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_0, ack => cp_elements(1766)); -- 
    -- CP-element group 1767 transition  output  bypass 
    -- predecessors 1764 
    -- successors 1768 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/cr
      -- 
    cp_elements(1767) <= cp_elements(1764);
    cr_15537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1767), ack => type_cast_2690_inst_req_1); -- 
    -- CP-element group 1768 transition  input  bypass 
    -- predecessors 1767 
    -- successors 1769 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/ca
      -- 
    ca_15538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_1, ack => cp_elements(1768)); -- 
    -- CP-element group 1769 join  transition  bypass 
    -- predecessors 1766 1768 
    -- successors 1774 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/$exit
      -- 
    cp_element_group_1769: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1769"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1766) & cp_elements(1768);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1769), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1770 fork  transition  bypass 
    -- predecessors 1763 
    -- successors 1771 1772 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/$entry
      -- 
    cp_elements(1770) <= cp_elements(1763);
    -- CP-element group 1771 transition  bypass 
    -- predecessors 1770 
    -- successors 1773 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/ra
      -- 
    cp_elements(1771) <= cp_elements(1770);
    -- CP-element group 1772 transition  bypass 
    -- predecessors 1770 
    -- successors 1773 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/ca
      -- 
    cp_elements(1772) <= cp_elements(1770);
    -- CP-element group 1773 join  transition  bypass 
    -- predecessors 1771 1772 
    -- successors 1774 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/$exit
      -- 
    cp_element_group_1773: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1773"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1771) & cp_elements(1772);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1773), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1774 join  transition  output  bypass 
    -- predecessors 1769 1773 
    -- successors 1775 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_req
      -- 
    cp_element_group_1774: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1774"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1769) & cp_elements(1773);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1774), clk => clk, reset => reset); --
    end block;
    phi_stmt_2687_req_15555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1774), ack => phi_stmt_2687_req_0); -- 
    -- CP-element group 1775 join  transition  bypass 
    -- predecessors 1762 1774 
    -- successors 1794 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1775: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1775"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1762) & cp_elements(1774);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1775), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1776 fork  transition  bypass 
    -- predecessors 38 
    -- successors 1777 1781 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1776) <= cp_elements(38);
    -- CP-element group 1777 fork  transition  bypass 
    -- predecessors 1776 
    -- successors 1778 1779 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/$entry
      -- 
    cp_elements(1777) <= cp_elements(1776);
    -- CP-element group 1778 transition  bypass 
    -- predecessors 1777 
    -- successors 1780 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Sample/ra
      -- 
    cp_elements(1778) <= cp_elements(1777);
    -- CP-element group 1779 transition  bypass 
    -- predecessors 1777 
    -- successors 1780 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/Update/ca
      -- 
    cp_elements(1779) <= cp_elements(1777);
    -- CP-element group 1780 join  transition  output  bypass 
    -- predecessors 1778 1779 
    -- successors 1793 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_sources/type_cast_2683/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2680/phi_stmt_2680_req
      -- 
    cp_element_group_1780: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1780"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1778) & cp_elements(1779);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1780), clk => clk, reset => reset); --
    end block;
    phi_stmt_2680_req_15581_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1780), ack => phi_stmt_2680_req_1); -- 
    -- CP-element group 1781 fork  transition  bypass 
    -- predecessors 1776 
    -- successors 1782 1786 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/$entry
      -- 
    cp_elements(1781) <= cp_elements(1776);
    -- CP-element group 1782 fork  transition  bypass 
    -- predecessors 1781 
    -- successors 1783 1784 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/$entry
      -- 
    cp_elements(1782) <= cp_elements(1781);
    -- CP-element group 1783 transition  bypass 
    -- predecessors 1782 
    -- successors 1785 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Sample/ra
      -- 
    cp_elements(1783) <= cp_elements(1782);
    -- CP-element group 1784 transition  bypass 
    -- predecessors 1782 
    -- successors 1785 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/Update/ca
      -- 
    cp_elements(1784) <= cp_elements(1782);
    -- CP-element group 1785 join  transition  bypass 
    -- predecessors 1783 1784 
    -- successors 1792 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2690/SplitProtocol/$exit
      -- 
    cp_element_group_1785: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1785"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1783) & cp_elements(1784);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1785), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1786 fork  transition  bypass 
    -- predecessors 1781 
    -- successors 1787 1789 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/$entry
      -- 
    cp_elements(1786) <= cp_elements(1781);
    -- CP-element group 1787 transition  output  bypass 
    -- predecessors 1786 
    -- successors 1788 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/rr
      -- 
    cp_elements(1787) <= cp_elements(1786);
    rr_15613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1787), ack => type_cast_2692_inst_req_0); -- 
    -- CP-element group 1788 transition  input  bypass 
    -- predecessors 1787 
    -- successors 1791 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Sample/ra
      -- 
    ra_15614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_0, ack => cp_elements(1788)); -- 
    -- CP-element group 1789 transition  output  bypass 
    -- predecessors 1786 
    -- successors 1790 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/cr
      -- 
    cp_elements(1789) <= cp_elements(1786);
    cr_15618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1789), ack => type_cast_2692_inst_req_1); -- 
    -- CP-element group 1790 transition  input  bypass 
    -- predecessors 1789 
    -- successors 1791 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/Update/ca
      -- 
    ca_15619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_1, ack => cp_elements(1790)); -- 
    -- CP-element group 1791 join  transition  bypass 
    -- predecessors 1788 1790 
    -- successors 1792 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/type_cast_2692/SplitProtocol/$exit
      -- 
    cp_element_group_1791: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1791"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1788) & cp_elements(1790);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1791), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1792 join  transition  output  bypass 
    -- predecessors 1785 1791 
    -- successors 1793 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/phi_stmt_2687/phi_stmt_2687_req
      -- 
    cp_element_group_1792: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1792"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1785) & cp_elements(1791);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1792), clk => clk, reset => reset); --
    end block;
    phi_stmt_2687_req_15620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1792), ack => phi_stmt_2687_req_1); -- 
    -- CP-element group 1793 join  transition  bypass 
    -- predecessors 1780 1792 
    -- successors 1794 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xix_xpreheader_udiv32x_xexitx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1793: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1793"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1780) & cp_elements(1792);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1793), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1794 merge  place  bypass 
    -- predecessors 1775 1793 
    -- successors 1795 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2679_PhiReqMerge
      -- 
    cp_elements(1794) <= OrReduce(cp_elements(1775) & cp_elements(1793));
    -- CP-element group 1795 fork  transition  bypass 
    -- predecessors 1794 
    -- successors 1796 1797 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2679_PhiAck/$entry
      -- 
    cp_elements(1795) <= cp_elements(1794);
    -- CP-element group 1796 transition  input  bypass 
    -- predecessors 1795 
    -- successors 1798 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2679_PhiAck/phi_stmt_2680_ack
      -- 
    phi_stmt_2680_ack_15625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2680_ack_0, ack => cp_elements(1796)); -- 
    -- CP-element group 1797 transition  input  bypass 
    -- predecessors 1795 
    -- successors 1798 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2679_PhiAck/phi_stmt_2687_ack
      -- 
    phi_stmt_2687_ack_15626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2687_ack_0, ack => cp_elements(1797)); -- 
    -- CP-element group 1798 join  transition  bypass 
    -- predecessors 1796 1797 
    -- successors 39 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2679_PhiAck/$exit
      -- 
    cp_element_group_1798: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1798"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1796) & cp_elements(1797);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1798), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1799 fork  transition  bypass 
    -- predecessors 725 
    -- successors 1800 1806 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1799) <= cp_elements(725);
    -- CP-element group 1800 fork  transition  bypass 
    -- predecessors 1799 
    -- successors 1801 1803 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/$entry
      -- 
    cp_elements(1800) <= cp_elements(1799);
    -- CP-element group 1801 transition  output  bypass 
    -- predecessors 1800 
    -- successors 1802 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Sample/rr
      -- 
    cp_elements(1801) <= cp_elements(1800);
    rr_15649_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1801), ack => type_cast_2741_inst_req_0); -- 
    -- CP-element group 1802 transition  input  bypass 
    -- predecessors 1801 
    -- successors 1805 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Sample/ra
      -- 
    ra_15650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2741_inst_ack_0, ack => cp_elements(1802)); -- 
    -- CP-element group 1803 transition  output  bypass 
    -- predecessors 1800 
    -- successors 1804 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Update/cr
      -- 
    cp_elements(1803) <= cp_elements(1800);
    cr_15654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1803), ack => type_cast_2741_inst_req_1); -- 
    -- CP-element group 1804 transition  input  bypass 
    -- predecessors 1803 
    -- successors 1805 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/Update/ca
      -- 
    ca_15655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2741_inst_ack_1, ack => cp_elements(1804)); -- 
    -- CP-element group 1805 join  transition  output  bypass 
    -- predecessors 1802 1804 
    -- successors 1812 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_sources/type_cast_2741/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2738/phi_stmt_2738_req
      -- 
    cp_element_group_1805: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1805"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1802) & cp_elements(1804);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1805), clk => clk, reset => reset); --
    end block;
    phi_stmt_2738_req_15656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1805), ack => phi_stmt_2738_req_0); -- 
    -- CP-element group 1806 fork  transition  bypass 
    -- predecessors 1799 
    -- successors 1807 1809 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/$entry
      -- 
    cp_elements(1806) <= cp_elements(1799);
    -- CP-element group 1807 transition  output  bypass 
    -- predecessors 1806 
    -- successors 1808 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Sample/rr
      -- 
    cp_elements(1807) <= cp_elements(1806);
    rr_15672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1807), ack => type_cast_2745_inst_req_0); -- 
    -- CP-element group 1808 transition  input  bypass 
    -- predecessors 1807 
    -- successors 1811 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Sample/ra
      -- 
    ra_15673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2745_inst_ack_0, ack => cp_elements(1808)); -- 
    -- CP-element group 1809 transition  output  bypass 
    -- predecessors 1806 
    -- successors 1810 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Update/cr
      -- 
    cp_elements(1809) <= cp_elements(1806);
    cr_15677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1809), ack => type_cast_2745_inst_req_1); -- 
    -- CP-element group 1810 transition  input  bypass 
    -- predecessors 1809 
    -- successors 1811 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/Update/ca
      -- 
    ca_15678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2745_inst_ack_1, ack => cp_elements(1810)); -- 
    -- CP-element group 1811 join  transition  output  bypass 
    -- predecessors 1808 1810 
    -- successors 1812 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_sources/type_cast_2745/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/phi_stmt_2742/phi_stmt_2742_req
      -- 
    cp_element_group_1811: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1811"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1808) & cp_elements(1810);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1811), clk => clk, reset => reset); --
    end block;
    phi_stmt_2742_req_15679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1811), ack => phi_stmt_2742_req_0); -- 
    -- CP-element group 1812 join  transition  bypass 
    -- predecessors 1805 1811 
    -- successors 1813 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1812: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1812"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1805) & cp_elements(1811);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1812), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1813 place  bypass 
    -- predecessors 1812 
    -- successors 1814 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2737_PhiReqMerge
      -- 
    cp_elements(1813) <= cp_elements(1812);
    -- CP-element group 1814 fork  transition  bypass 
    -- predecessors 1813 
    -- successors 1815 1816 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2737_PhiAck/$entry
      -- 
    cp_elements(1814) <= cp_elements(1813);
    -- CP-element group 1815 transition  input  bypass 
    -- predecessors 1814 
    -- successors 1817 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2737_PhiAck/phi_stmt_2738_ack
      -- 
    phi_stmt_2738_ack_15684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2738_ack_0, ack => cp_elements(1815)); -- 
    -- CP-element group 1816 transition  input  bypass 
    -- predecessors 1814 
    -- successors 1817 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2737_PhiAck/phi_stmt_2742_ack
      -- 
    phi_stmt_2742_ack_15685_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2742_ack_0, ack => cp_elements(1816)); -- 
    -- CP-element group 1817 join  transition  bypass 
    -- predecessors 1815 1816 
    -- successors 41 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2737_PhiAck/$exit
      -- 
    cp_element_group_1817: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1817"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1815) & cp_elements(1816);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1817), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1818 fork  transition  bypass 
    -- predecessors 691 
    -- successors 1819 1831 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1818) <= cp_elements(691);
    -- CP-element group 1819 fork  transition  bypass 
    -- predecessors 1818 
    -- successors 1820 1824 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/$entry
      -- 
    cp_elements(1819) <= cp_elements(1818);
    -- CP-element group 1820 fork  transition  bypass 
    -- predecessors 1819 
    -- successors 1821 1822 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/$entry
      -- 
    cp_elements(1820) <= cp_elements(1819);
    -- CP-element group 1821 transition  bypass 
    -- predecessors 1820 
    -- successors 1823 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/ra
      -- 
    cp_elements(1821) <= cp_elements(1820);
    -- CP-element group 1822 transition  bypass 
    -- predecessors 1820 
    -- successors 1823 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/ca
      -- 
    cp_elements(1822) <= cp_elements(1820);
    -- CP-element group 1823 join  transition  bypass 
    -- predecessors 1821 1822 
    -- successors 1830 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/$exit
      -- 
    cp_element_group_1823: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1823"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1821) & cp_elements(1822);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1823), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1824 fork  transition  bypass 
    -- predecessors 1819 
    -- successors 1825 1827 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/$entry
      -- 
    cp_elements(1824) <= cp_elements(1819);
    -- CP-element group 1825 transition  output  bypass 
    -- predecessors 1824 
    -- successors 1826 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/rr
      -- 
    cp_elements(1825) <= cp_elements(1824);
    rr_15720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1825), ack => type_cast_2776_inst_req_0); -- 
    -- CP-element group 1826 transition  input  bypass 
    -- predecessors 1825 
    -- successors 1829 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/ra
      -- 
    ra_15721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_0, ack => cp_elements(1826)); -- 
    -- CP-element group 1827 transition  output  bypass 
    -- predecessors 1824 
    -- successors 1828 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/cr
      -- 
    cp_elements(1827) <= cp_elements(1824);
    cr_15725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1827), ack => type_cast_2776_inst_req_1); -- 
    -- CP-element group 1828 transition  input  bypass 
    -- predecessors 1827 
    -- successors 1829 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/ca
      -- 
    ca_15726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_1, ack => cp_elements(1828)); -- 
    -- CP-element group 1829 join  transition  bypass 
    -- predecessors 1826 1828 
    -- successors 1830 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/$exit
      -- 
    cp_element_group_1829: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1829"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1826) & cp_elements(1828);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1829), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1830 join  transition  output  bypass 
    -- predecessors 1823 1829 
    -- successors 1843 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_req
      -- 
    cp_element_group_1830: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1830"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1823) & cp_elements(1829);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1830), clk => clk, reset => reset); --
    end block;
    phi_stmt_2771_req_15727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1830), ack => phi_stmt_2771_req_1); -- 
    -- CP-element group 1831 fork  transition  bypass 
    -- predecessors 1818 
    -- successors 1832 1836 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/$entry
      -- 
    cp_elements(1831) <= cp_elements(1818);
    -- CP-element group 1832 fork  transition  bypass 
    -- predecessors 1831 
    -- successors 1833 1834 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/$entry
      -- 
    cp_elements(1832) <= cp_elements(1831);
    -- CP-element group 1833 transition  bypass 
    -- predecessors 1832 
    -- successors 1835 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/ra
      -- 
    cp_elements(1833) <= cp_elements(1832);
    -- CP-element group 1834 transition  bypass 
    -- predecessors 1832 
    -- successors 1835 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/ca
      -- 
    cp_elements(1834) <= cp_elements(1832);
    -- CP-element group 1835 join  transition  bypass 
    -- predecessors 1833 1834 
    -- successors 1842 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/$exit
      -- 
    cp_element_group_1835: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1835"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1833) & cp_elements(1834);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1835), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1836 fork  transition  bypass 
    -- predecessors 1831 
    -- successors 1837 1839 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/$entry
      -- 
    cp_elements(1836) <= cp_elements(1831);
    -- CP-element group 1837 transition  output  bypass 
    -- predecessors 1836 
    -- successors 1838 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/rr
      -- 
    cp_elements(1837) <= cp_elements(1836);
    rr_15759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1837), ack => type_cast_2782_inst_req_0); -- 
    -- CP-element group 1838 transition  input  bypass 
    -- predecessors 1837 
    -- successors 1841 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/ra
      -- 
    ra_15760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_0, ack => cp_elements(1838)); -- 
    -- CP-element group 1839 transition  output  bypass 
    -- predecessors 1836 
    -- successors 1840 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/cr
      -- 
    cp_elements(1839) <= cp_elements(1836);
    cr_15764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1839), ack => type_cast_2782_inst_req_1); -- 
    -- CP-element group 1840 transition  input  bypass 
    -- predecessors 1839 
    -- successors 1841 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/ca
      -- 
    ca_15765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_1, ack => cp_elements(1840)); -- 
    -- CP-element group 1841 join  transition  bypass 
    -- predecessors 1838 1840 
    -- successors 1842 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/$exit
      -- 
    cp_element_group_1841: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1841"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1838) & cp_elements(1840);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1841), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1842 join  transition  output  bypass 
    -- predecessors 1835 1841 
    -- successors 1843 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_req
      -- 
    cp_element_group_1842: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1842"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1835) & cp_elements(1841);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1842), clk => clk, reset => reset); --
    end block;
    phi_stmt_2777_req_15766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1842), ack => phi_stmt_2777_req_1); -- 
    -- CP-element group 1843 join  transition  bypass 
    -- predecessors 1830 1842 
    -- successors 1870 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1843: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1843"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1830) & cp_elements(1842);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1844 fork  transition  bypass 
    -- predecessors 743 
    -- successors 1845 1857 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1844) <= cp_elements(743);
    -- CP-element group 1845 fork  transition  bypass 
    -- predecessors 1844 
    -- successors 1846 1852 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/$entry
      -- 
    cp_elements(1845) <= cp_elements(1844);
    -- CP-element group 1846 fork  transition  bypass 
    -- predecessors 1845 
    -- successors 1847 1849 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/$entry
      -- 
    cp_elements(1846) <= cp_elements(1845);
    -- CP-element group 1847 transition  output  bypass 
    -- predecessors 1846 
    -- successors 1848 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1847) <= cp_elements(1846);
    rr_15785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1847), ack => type_cast_2774_inst_req_0); -- 
    -- CP-element group 1848 transition  input  bypass 
    -- predecessors 1847 
    -- successors 1851 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Sample/$exit
      -- 
    ra_15786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2774_inst_ack_0, ack => cp_elements(1848)); -- 
    -- CP-element group 1849 transition  output  bypass 
    -- predecessors 1846 
    -- successors 1850 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/$entry
      -- 
    cp_elements(1849) <= cp_elements(1846);
    cr_15790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1849), ack => type_cast_2774_inst_req_1); -- 
    -- CP-element group 1850 transition  input  bypass 
    -- predecessors 1849 
    -- successors 1851 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/Update/$exit
      -- 
    ca_15791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2774_inst_ack_1, ack => cp_elements(1850)); -- 
    -- CP-element group 1851 join  transition  bypass 
    -- predecessors 1848 1850 
    -- successors 1856 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2774/$exit
      -- 
    cp_element_group_1851: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1851"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1848) & cp_elements(1850);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1851), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1852 fork  transition  bypass 
    -- predecessors 1845 
    -- successors 1853 1854 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/$entry
      -- 
    cp_elements(1852) <= cp_elements(1845);
    -- CP-element group 1853 transition  bypass 
    -- predecessors 1852 
    -- successors 1855 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Sample/ra
      -- 
    cp_elements(1853) <= cp_elements(1852);
    -- CP-element group 1854 transition  bypass 
    -- predecessors 1852 
    -- successors 1855 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/Update/ca
      -- 
    cp_elements(1854) <= cp_elements(1852);
    -- CP-element group 1855 join  transition  bypass 
    -- predecessors 1853 1854 
    -- successors 1856 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/type_cast_2776/$exit
      -- 
    cp_element_group_1855: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1855"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1853) & cp_elements(1854);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1855), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1856 join  transition  output  bypass 
    -- predecessors 1851 1855 
    -- successors 1869 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2771/phi_stmt_2771_req
      -- 
    cp_element_group_1856: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1856"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1851) & cp_elements(1855);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1856), clk => clk, reset => reset); --
    end block;
    phi_stmt_2771_req_15808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1856), ack => phi_stmt_2771_req_0); -- 
    -- CP-element group 1857 fork  transition  bypass 
    -- predecessors 1844 
    -- successors 1858 1864 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/$entry
      -- 
    cp_elements(1857) <= cp_elements(1844);
    -- CP-element group 1858 fork  transition  bypass 
    -- predecessors 1857 
    -- successors 1859 1861 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/$entry
      -- 
    cp_elements(1858) <= cp_elements(1857);
    -- CP-element group 1859 transition  output  bypass 
    -- predecessors 1858 
    -- successors 1860 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1859) <= cp_elements(1858);
    rr_15824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1859), ack => type_cast_2780_inst_req_0); -- 
    -- CP-element group 1860 transition  input  bypass 
    -- predecessors 1859 
    -- successors 1863 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Sample/$exit
      -- 
    ra_15825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_0, ack => cp_elements(1860)); -- 
    -- CP-element group 1861 transition  output  bypass 
    -- predecessors 1858 
    -- successors 1862 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/$entry
      -- 
    cp_elements(1861) <= cp_elements(1858);
    cr_15829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1861), ack => type_cast_2780_inst_req_1); -- 
    -- CP-element group 1862 transition  input  bypass 
    -- predecessors 1861 
    -- successors 1863 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/Update/$exit
      -- 
    ca_15830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_1, ack => cp_elements(1862)); -- 
    -- CP-element group 1863 join  transition  bypass 
    -- predecessors 1860 1862 
    -- successors 1868 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2780/$exit
      -- 
    cp_element_group_1863: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1863"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1860) & cp_elements(1862);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1863), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1864 fork  transition  bypass 
    -- predecessors 1857 
    -- successors 1865 1866 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/$entry
      -- 
    cp_elements(1864) <= cp_elements(1857);
    -- CP-element group 1865 transition  bypass 
    -- predecessors 1864 
    -- successors 1867 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1865) <= cp_elements(1864);
    -- CP-element group 1866 transition  bypass 
    -- predecessors 1864 
    -- successors 1867 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/Update/$entry
      -- 
    cp_elements(1866) <= cp_elements(1864);
    -- CP-element group 1867 join  transition  bypass 
    -- predecessors 1865 1866 
    -- successors 1868 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/type_cast_2782/$exit
      -- 
    cp_element_group_1867: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1867"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1865) & cp_elements(1866);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1867), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1868 join  transition  output  bypass 
    -- predecessors 1863 1867 
    -- successors 1869 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_req
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/phi_stmt_2777_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/phi_stmt_2777/$exit
      -- 
    cp_element_group_1868: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1868"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1863) & cp_elements(1867);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1868), clk => clk, reset => reset); --
    end block;
    phi_stmt_2777_req_15847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1868), ack => phi_stmt_2777_req_0); -- 
    -- CP-element group 1869 join  transition  bypass 
    -- predecessors 1856 1868 
    -- successors 1870 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xix_xi_xx_xcritedgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1869: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1869"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1856) & cp_elements(1868);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1869), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1870 merge  place  bypass 
    -- predecessors 1843 1869 
    -- successors 1871 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2770_PhiReqMerge
      -- 
    cp_elements(1870) <= OrReduce(cp_elements(1843) & cp_elements(1869));
    -- CP-element group 1871 fork  transition  bypass 
    -- predecessors 1870 
    -- successors 1872 1873 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2770_PhiAck/$entry
      -- 
    cp_elements(1871) <= cp_elements(1870);
    -- CP-element group 1872 transition  input  bypass 
    -- predecessors 1871 
    -- successors 1874 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2770_PhiAck/phi_stmt_2771_ack
      -- 
    phi_stmt_2771_ack_15852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2771_ack_0, ack => cp_elements(1872)); -- 
    -- CP-element group 1873 transition  input  bypass 
    -- predecessors 1871 
    -- successors 1874 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2770_PhiAck/phi_stmt_2777_ack
      -- 
    phi_stmt_2777_ack_15853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2777_ack_0, ack => cp_elements(1873)); -- 
    -- CP-element group 1874 join  transition  bypass 
    -- predecessors 1872 1873 
    -- successors 42 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2770_PhiAck/$exit
      -- 
    cp_element_group_1874: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1874"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1872) & cp_elements(1873);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1874), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1875 transition  bypass 
    -- predecessors 527 
    -- successors 1877 
    -- members (4) 
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/$entry
      -- 
    cp_elements(1875) <= cp_elements(527);
    -- CP-element group 1876 transition  bypass 
    -- predecessors 527 
    -- successors 1877 
    -- members (4) 
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/$entry
      -- 
    cp_elements(1876) <= cp_elements(527);
    -- CP-element group 1877 join  transition  output  bypass 
    -- predecessors 1875 1876 
    -- successors 1883 
    -- members (6) 
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_req
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/$exit
      -- 	branch_block_stmt_1659/omega_calcx_xexit_iq_err_calcx_xexit_PhiReq/$exit
      -- 
    cp_element_group_1877: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1877"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1875) & cp_elements(1876);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1877), clk => clk, reset => reset); --
    end block;
    phi_stmt_2818_req_15879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1877), ack => phi_stmt_2818_req_1); -- 
    -- CP-element group 1878 transition  output  bypass 
    -- predecessors 767 
    -- successors 1879 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/rr
      -- 
    cp_elements(1878) <= cp_elements(767);
    rr_15898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1878), ack => type_cast_2821_inst_req_0); -- 
    -- CP-element group 1879 transition  input  bypass 
    -- predecessors 1878 
    -- successors 1882 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/ra
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Sample/$exit
      -- 
    ra_15899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2821_inst_ack_0, ack => cp_elements(1879)); -- 
    -- CP-element group 1880 transition  output  bypass 
    -- predecessors 767 
    -- successors 1881 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/$entry
      -- 
    cp_elements(1880) <= cp_elements(767);
    cr_15903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1880), ack => type_cast_2821_inst_req_1); -- 
    -- CP-element group 1881 transition  input  bypass 
    -- predecessors 1880 
    -- successors 1882 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/ca
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/Update/$exit
      -- 
    ca_15904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2821_inst_ack_1, ack => cp_elements(1881)); -- 
    -- CP-element group 1882 join  transition  output  bypass 
    -- predecessors 1879 1881 
    -- successors 1883 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_req
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/type_cast_2821/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/phi_stmt_2818_sources/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/phi_stmt_2818/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xix_xi_iq_err_calcx_xexit_PhiReq/$exit
      -- 
    cp_element_group_1882: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1882"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1879) & cp_elements(1881);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1882), clk => clk, reset => reset); --
    end block;
    phi_stmt_2818_req_15905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1882), ack => phi_stmt_2818_req_0); -- 
    -- CP-element group 1883 merge  place  bypass 
    -- predecessors 1877 1882 
    -- successors 1884 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2817_PhiReqMerge
      -- 
    cp_elements(1883) <= OrReduce(cp_elements(1877) & cp_elements(1882));
    -- CP-element group 1884 transition  bypass 
    -- predecessors 1883 
    -- successors 1885 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2817_PhiAck/$entry
      -- 
    cp_elements(1884) <= cp_elements(1883);
    -- CP-element group 1885 transition  place  input  bypass 
    -- predecessors 1884 
    -- successors 768 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2831_to_assign_stmt_2865__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2817__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2817_PhiAck/phi_stmt_2818_ack
      -- 	branch_block_stmt_1659/merge_stmt_2817_PhiAck/$exit
      -- 
    phi_stmt_2818_ack_15910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2818_ack_0, ack => cp_elements(1885)); -- 
    -- CP-element group 1886 transition  bypass 
    -- predecessors 811 
    -- successors 1888 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/ra
      -- 
    cp_elements(1886) <= cp_elements(811);
    -- CP-element group 1887 transition  bypass 
    -- predecessors 811 
    -- successors 1888 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/ca
      -- 
    cp_elements(1887) <= cp_elements(811);
    -- CP-element group 1888 join  transition  output  bypass 
    -- predecessors 1886 1887 
    -- successors 1897 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_42_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_req
      -- 
    cp_element_group_1888: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1888"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1886) & cp_elements(1887);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1888), clk => clk, reset => reset); --
    end block;
    phi_stmt_2888_req_15960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1888), ack => phi_stmt_2888_req_2); -- 
    -- CP-element group 1889 transition  output  bypass 
    -- predecessors 44 
    -- successors 1890 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/rr
      -- 
    cp_elements(1889) <= cp_elements(44);
    rr_15979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1889), ack => type_cast_2891_inst_req_0); -- 
    -- CP-element group 1890 transition  input  bypass 
    -- predecessors 1889 
    -- successors 1893 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/ra
      -- 
    ra_15980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2891_inst_ack_0, ack => cp_elements(1890)); -- 
    -- CP-element group 1891 transition  output  bypass 
    -- predecessors 44 
    -- successors 1892 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/cr
      -- 
    cp_elements(1891) <= cp_elements(44);
    cr_15984_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1891), ack => type_cast_2891_inst_req_1); -- 
    -- CP-element group 1892 transition  input  bypass 
    -- predecessors 1891 
    -- successors 1893 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/ca
      -- 
    ca_15985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2891_inst_ack_1, ack => cp_elements(1892)); -- 
    -- CP-element group 1893 join  transition  output  bypass 
    -- predecessors 1890 1892 
    -- successors 1897 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_43_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_req
      -- 
    cp_element_group_1893: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1893"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1890) & cp_elements(1892);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1893), clk => clk, reset => reset); --
    end block;
    phi_stmt_2888_req_15986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1893), ack => phi_stmt_2888_req_0); -- 
    -- CP-element group 1894 transition  bypass 
    -- predecessors 799 
    -- successors 1896 
    -- members (4) 
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Sample/ra
      -- 
    cp_elements(1894) <= cp_elements(799);
    -- CP-element group 1895 transition  bypass 
    -- predecessors 799 
    -- successors 1896 
    -- members (4) 
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/Update/ca
      -- 
    cp_elements(1895) <= cp_elements(799);
    -- CP-element group 1896 join  transition  output  bypass 
    -- predecessors 1894 1895 
    -- successors 1897 
    -- members (6) 
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_sources/type_cast_2891/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/iq_err_calcx_xexit_bb_44_PhiReq/phi_stmt_2888/phi_stmt_2888_req
      -- 
    cp_element_group_1896: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1896"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1894) & cp_elements(1895);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1896), clk => clk, reset => reset); --
    end block;
    phi_stmt_2888_req_16012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1896), ack => phi_stmt_2888_req_1); -- 
    -- CP-element group 1897 merge  place  bypass 
    -- predecessors 1888 1893 1896 
    -- successors 1898 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2887_PhiReqMerge
      -- 
    cp_elements(1897) <= OrReduce(cp_elements(1888) & cp_elements(1893) & cp_elements(1896));
    -- CP-element group 1898 transition  bypass 
    -- predecessors 1897 
    -- successors 1899 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2887_PhiAck/$entry
      -- 
    cp_elements(1898) <= cp_elements(1897);
    -- CP-element group 1899 transition  place  input  bypass 
    -- predecessors 1898 
    -- successors 814 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_2904_to_assign_stmt_2915__entry__
      -- 	branch_block_stmt_1659/merge_stmt_2887__exit__
      -- 	branch_block_stmt_1659/merge_stmt_2887_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2887_PhiAck/phi_stmt_2888_ack
      -- 
    phi_stmt_2888_ack_16017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2888_ack_0, ack => cp_elements(1899)); -- 
    -- CP-element group 1900 transition  bypass 
    -- predecessors 831 
    -- successors 1902 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/ra
      -- 
    cp_elements(1900) <= cp_elements(831);
    -- CP-element group 1901 transition  bypass 
    -- predecessors 831 
    -- successors 1902 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/ca
      -- 
    cp_elements(1901) <= cp_elements(831);
    -- CP-element group 1902 join  transition  output  bypass 
    -- predecessors 1900 1901 
    -- successors 1911 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_44_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_req
      -- 
    cp_element_group_1902: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1902"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1900) & cp_elements(1901);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1902), clk => clk, reset => reset); --
    end block;
    phi_stmt_2949_req_16071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1902), ack => phi_stmt_2949_req_1); -- 
    -- CP-element group 1903 transition  bypass 
    -- predecessors 843 
    -- successors 1905 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/ra
      -- 
    cp_elements(1903) <= cp_elements(843);
    -- CP-element group 1904 transition  bypass 
    -- predecessors 843 
    -- successors 1905 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/ca
      -- 
    cp_elements(1904) <= cp_elements(843);
    -- CP-element group 1905 join  transition  output  bypass 
    -- predecessors 1903 1904 
    -- successors 1911 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_45_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_req
      -- 
    cp_element_group_1905: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1905"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1903) & cp_elements(1904);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1905), clk => clk, reset => reset); --
    end block;
    phi_stmt_2949_req_16097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1905), ack => phi_stmt_2949_req_2); -- 
    -- CP-element group 1906 transition  output  bypass 
    -- predecessors 857 
    -- successors 1907 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/rr
      -- 
    cp_elements(1906) <= cp_elements(857);
    rr_16116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1906), ack => type_cast_2952_inst_req_0); -- 
    -- CP-element group 1907 transition  input  bypass 
    -- predecessors 1906 
    -- successors 1910 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Sample/ra
      -- 
    ra_16117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2952_inst_ack_0, ack => cp_elements(1907)); -- 
    -- CP-element group 1908 transition  output  bypass 
    -- predecessors 857 
    -- successors 1909 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/cr
      -- 
    cp_elements(1908) <= cp_elements(857);
    cr_16121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1908), ack => type_cast_2952_inst_req_1); -- 
    -- CP-element group 1909 transition  input  bypass 
    -- predecessors 1908 
    -- successors 1910 
    -- members (2) 
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/Update/ca
      -- 
    ca_16122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2952_inst_ack_1, ack => cp_elements(1909)); -- 
    -- CP-element group 1910 join  transition  output  bypass 
    -- predecessors 1907 1909 
    -- successors 1911 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_sources/type_cast_2952/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_46_xx_xthread_PhiReq/phi_stmt_2949/phi_stmt_2949_req
      -- 
    cp_element_group_1910: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1910"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1907) & cp_elements(1909);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1910), clk => clk, reset => reset); --
    end block;
    phi_stmt_2949_req_16123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1910), ack => phi_stmt_2949_req_0); -- 
    -- CP-element group 1911 merge  place  bypass 
    -- predecessors 1902 1905 1910 
    -- successors 1912 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2948_PhiReqMerge
      -- 
    cp_elements(1911) <= OrReduce(cp_elements(1902) & cp_elements(1905) & cp_elements(1910));
    -- CP-element group 1912 transition  bypass 
    -- predecessors 1911 
    -- successors 1913 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2948_PhiAck/$entry
      -- 
    cp_elements(1912) <= cp_elements(1911);
    -- CP-element group 1913 transition  input  bypass 
    -- predecessors 1912 
    -- successors 47 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_2948_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_2948_PhiAck/phi_stmt_2949_ack
      -- 
    phi_stmt_2949_ack_16128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2949_ack_0, ack => cp_elements(1913)); -- 
    -- CP-element group 1914 fork  transition  bypass 
    -- predecessors 932 
    -- successors 1915 1927 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1914) <= cp_elements(932);
    -- CP-element group 1915 fork  transition  bypass 
    -- predecessors 1914 
    -- successors 1916 1922 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/$entry
      -- 
    cp_elements(1915) <= cp_elements(1914);
    -- CP-element group 1916 fork  transition  bypass 
    -- predecessors 1915 
    -- successors 1917 1919 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/$entry
      -- 
    cp_elements(1916) <= cp_elements(1915);
    -- CP-element group 1917 transition  output  bypass 
    -- predecessors 1916 
    -- successors 1918 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/rr
      -- 
    cp_elements(1917) <= cp_elements(1916);
    rr_16147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1917), ack => type_cast_2987_inst_req_0); -- 
    -- CP-element group 1918 transition  input  bypass 
    -- predecessors 1917 
    -- successors 1921 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/ra
      -- 
    ra_16148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2987_inst_ack_0, ack => cp_elements(1918)); -- 
    -- CP-element group 1919 transition  output  bypass 
    -- predecessors 1916 
    -- successors 1920 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/cr
      -- 
    cp_elements(1919) <= cp_elements(1916);
    cr_16152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1919), ack => type_cast_2987_inst_req_1); -- 
    -- CP-element group 1920 transition  input  bypass 
    -- predecessors 1919 
    -- successors 1921 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/ca
      -- 
    ca_16153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2987_inst_ack_1, ack => cp_elements(1920)); -- 
    -- CP-element group 1921 join  transition  bypass 
    -- predecessors 1918 1920 
    -- successors 1926 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/$exit
      -- 
    cp_element_group_1921: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1921"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1918) & cp_elements(1920);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1921), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1922 fork  transition  bypass 
    -- predecessors 1915 
    -- successors 1923 1924 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/$entry
      -- 
    cp_elements(1922) <= cp_elements(1915);
    -- CP-element group 1923 transition  bypass 
    -- predecessors 1922 
    -- successors 1925 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/ra
      -- 
    cp_elements(1923) <= cp_elements(1922);
    -- CP-element group 1924 transition  bypass 
    -- predecessors 1922 
    -- successors 1925 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/ca
      -- 
    cp_elements(1924) <= cp_elements(1922);
    -- CP-element group 1925 join  transition  bypass 
    -- predecessors 1923 1924 
    -- successors 1926 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/$exit
      -- 
    cp_element_group_1925: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1925"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1923) & cp_elements(1924);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1926 join  transition  output  bypass 
    -- predecessors 1921 1925 
    -- successors 1933 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_req
      -- 
    cp_element_group_1926: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1926"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1921) & cp_elements(1925);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1926), clk => clk, reset => reset); --
    end block;
    phi_stmt_2984_req_16170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1926), ack => phi_stmt_2984_req_0); -- 
    -- CP-element group 1927 fork  transition  bypass 
    -- predecessors 1914 
    -- successors 1928 1930 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$entry
      -- 
    cp_elements(1927) <= cp_elements(1914);
    -- CP-element group 1928 transition  output  bypass 
    -- predecessors 1927 
    -- successors 1929 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/rr
      -- 
    cp_elements(1928) <= cp_elements(1927);
    rr_16186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1928), ack => type_cast_2993_inst_req_0); -- 
    -- CP-element group 1929 transition  input  bypass 
    -- predecessors 1928 
    -- successors 1932 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/ra
      -- 
    ra_16187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_0, ack => cp_elements(1929)); -- 
    -- CP-element group 1930 transition  output  bypass 
    -- predecessors 1927 
    -- successors 1931 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/cr
      -- 
    cp_elements(1930) <= cp_elements(1927);
    cr_16191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1930), ack => type_cast_2993_inst_req_1); -- 
    -- CP-element group 1931 transition  input  bypass 
    -- predecessors 1930 
    -- successors 1932 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/ca
      -- 
    ca_16192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2993_inst_ack_1, ack => cp_elements(1931)); -- 
    -- CP-element group 1932 join  transition  output  bypass 
    -- predecessors 1929 1931 
    -- successors 1933 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- 
    cp_element_group_1932: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1932"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1929) & cp_elements(1931);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1932), clk => clk, reset => reset); --
    end block;
    phi_stmt_2990_req_16193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1932), ack => phi_stmt_2990_req_0); -- 
    -- CP-element group 1933 join  transition  bypass 
    -- predecessors 1926 1932 
    -- successors 1952 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_bbx_xnph7x_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1933: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1933"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1926) & cp_elements(1932);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1933), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1934 fork  transition  bypass 
    -- predecessors 871 
    -- successors 1935 1947 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1934) <= cp_elements(871);
    -- CP-element group 1935 fork  transition  bypass 
    -- predecessors 1934 
    -- successors 1936 1940 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/$entry
      -- 
    cp_elements(1935) <= cp_elements(1934);
    -- CP-element group 1936 fork  transition  bypass 
    -- predecessors 1935 
    -- successors 1937 1938 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/$entry
      -- 
    cp_elements(1936) <= cp_elements(1935);
    -- CP-element group 1937 transition  bypass 
    -- predecessors 1936 
    -- successors 1939 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Sample/ra
      -- 
    cp_elements(1937) <= cp_elements(1936);
    -- CP-element group 1938 transition  bypass 
    -- predecessors 1936 
    -- successors 1939 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/Update/ca
      -- 
    cp_elements(1938) <= cp_elements(1936);
    -- CP-element group 1939 join  transition  bypass 
    -- predecessors 1937 1938 
    -- successors 1946 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2987/SplitProtocol/$exit
      -- 
    cp_element_group_1939: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1939"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1937) & cp_elements(1938);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1939), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1940 fork  transition  bypass 
    -- predecessors 1935 
    -- successors 1941 1943 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/$entry
      -- 
    cp_elements(1940) <= cp_elements(1935);
    -- CP-element group 1941 transition  output  bypass 
    -- predecessors 1940 
    -- successors 1942 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/rr
      -- 
    cp_elements(1941) <= cp_elements(1940);
    rr_16228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1941), ack => type_cast_2989_inst_req_0); -- 
    -- CP-element group 1942 transition  input  bypass 
    -- predecessors 1941 
    -- successors 1945 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Sample/ra
      -- 
    ra_16229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2989_inst_ack_0, ack => cp_elements(1942)); -- 
    -- CP-element group 1943 transition  output  bypass 
    -- predecessors 1940 
    -- successors 1944 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/cr
      -- 
    cp_elements(1943) <= cp_elements(1940);
    cr_16233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1943), ack => type_cast_2989_inst_req_1); -- 
    -- CP-element group 1944 transition  input  bypass 
    -- predecessors 1943 
    -- successors 1945 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/Update/ca
      -- 
    ca_16234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2989_inst_ack_1, ack => cp_elements(1944)); -- 
    -- CP-element group 1945 join  transition  bypass 
    -- predecessors 1942 1944 
    -- successors 1946 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/type_cast_2989/SplitProtocol/$exit
      -- 
    cp_element_group_1945: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1945"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1942) & cp_elements(1944);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1945), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1946 join  transition  output  bypass 
    -- predecessors 1939 1945 
    -- successors 1951 
    -- members (3) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_sources/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2984/phi_stmt_2984_req
      -- 
    cp_element_group_1946: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1946"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1939) & cp_elements(1945);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1946), clk => clk, reset => reset); --
    end block;
    phi_stmt_2984_req_16235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1946), ack => phi_stmt_2984_req_1); -- 
    -- CP-element group 1947 fork  transition  bypass 
    -- predecessors 1934 
    -- successors 1948 1949 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$entry
      -- 
    cp_elements(1947) <= cp_elements(1934);
    -- CP-element group 1948 transition  bypass 
    -- predecessors 1947 
    -- successors 1950 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Sample/ra
      -- 
    cp_elements(1948) <= cp_elements(1947);
    -- CP-element group 1949 transition  bypass 
    -- predecessors 1947 
    -- successors 1950 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/Update/ca
      -- 
    cp_elements(1949) <= cp_elements(1947);
    -- CP-element group 1950 join  transition  output  bypass 
    -- predecessors 1948 1949 
    -- successors 1951 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_sources/type_cast_2993/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/phi_stmt_2990/phi_stmt_2990_req
      -- 
    cp_element_group_1950: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1950"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1948) & cp_elements(1949);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1950), clk => clk, reset => reset); --
    end block;
    phi_stmt_2990_req_16258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1950), ack => phi_stmt_2990_req_1); -- 
    -- CP-element group 1951 join  transition  bypass 
    -- predecessors 1946 1950 
    -- successors 1952 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_xthread_bbx_xnph7x_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1951: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1951"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1946) & cp_elements(1950);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1951), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1952 merge  place  bypass 
    -- predecessors 1933 1951 
    -- successors 1953 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2983_PhiReqMerge
      -- 
    cp_elements(1952) <= OrReduce(cp_elements(1933) & cp_elements(1951));
    -- CP-element group 1953 fork  transition  bypass 
    -- predecessors 1952 
    -- successors 1954 1955 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2983_PhiAck/$entry
      -- 
    cp_elements(1953) <= cp_elements(1952);
    -- CP-element group 1954 transition  input  bypass 
    -- predecessors 1953 
    -- successors 1956 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2983_PhiAck/phi_stmt_2984_ack
      -- 
    phi_stmt_2984_ack_16263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2984_ack_0, ack => cp_elements(1954)); -- 
    -- CP-element group 1955 transition  input  bypass 
    -- predecessors 1953 
    -- successors 1956 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2983_PhiAck/phi_stmt_2990_ack
      -- 
    phi_stmt_2990_ack_16264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2990_ack_0, ack => cp_elements(1955)); -- 
    -- CP-element group 1956 join  transition  bypass 
    -- predecessors 1954 1955 
    -- successors 48 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_2983_PhiAck/$exit
      -- 
    cp_element_group_1956: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1956"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1954) & cp_elements(1955);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1956), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1957 fork  transition  bypass 
    -- predecessors 906 
    -- successors 1958 1964 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1957) <= cp_elements(906);
    -- CP-element group 1958 fork  transition  bypass 
    -- predecessors 1957 
    -- successors 1959 1961 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/$entry
      -- 
    cp_elements(1958) <= cp_elements(1957);
    -- CP-element group 1959 transition  output  bypass 
    -- predecessors 1958 
    -- successors 1960 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/rr
      -- 
    cp_elements(1959) <= cp_elements(1958);
    rr_16295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1959), ack => type_cast_3022_inst_req_0); -- 
    -- CP-element group 1960 transition  input  bypass 
    -- predecessors 1959 
    -- successors 1963 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/ra
      -- 
    ra_16296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3022_inst_ack_0, ack => cp_elements(1960)); -- 
    -- CP-element group 1961 transition  output  bypass 
    -- predecessors 1958 
    -- successors 1962 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/cr
      -- 
    cp_elements(1961) <= cp_elements(1958);
    cr_16300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1961), ack => type_cast_3022_inst_req_1); -- 
    -- CP-element group 1962 transition  input  bypass 
    -- predecessors 1961 
    -- successors 1963 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/ca
      -- 
    ca_16301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3022_inst_ack_1, ack => cp_elements(1962)); -- 
    -- CP-element group 1963 join  transition  output  bypass 
    -- predecessors 1960 1962 
    -- successors 1970 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_req
      -- 
    cp_element_group_1963: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1963"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1960) & cp_elements(1962);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1963), clk => clk, reset => reset); --
    end block;
    phi_stmt_3019_req_16302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1963), ack => phi_stmt_3019_req_0); -- 
    -- CP-element group 1964 fork  transition  bypass 
    -- predecessors 1957 
    -- successors 1965 1967 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/$entry
      -- 
    cp_elements(1964) <= cp_elements(1957);
    -- CP-element group 1965 transition  output  bypass 
    -- predecessors 1964 
    -- successors 1966 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/rr
      -- 
    cp_elements(1965) <= cp_elements(1964);
    rr_16318_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1965), ack => type_cast_3029_inst_req_0); -- 
    -- CP-element group 1966 transition  input  bypass 
    -- predecessors 1965 
    -- successors 1969 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/ra
      -- 
    ra_16319_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3029_inst_ack_0, ack => cp_elements(1966)); -- 
    -- CP-element group 1967 transition  output  bypass 
    -- predecessors 1964 
    -- successors 1968 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/cr
      -- 
    cp_elements(1967) <= cp_elements(1964);
    cr_16323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1967), ack => type_cast_3029_inst_req_1); -- 
    -- CP-element group 1968 transition  input  bypass 
    -- predecessors 1967 
    -- successors 1969 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/ca
      -- 
    ca_16324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3029_inst_ack_1, ack => cp_elements(1968)); -- 
    -- CP-element group 1969 join  transition  output  bypass 
    -- predecessors 1966 1968 
    -- successors 1970 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_req
      -- 
    cp_element_group_1969: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1969"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1966) & cp_elements(1968);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1969), clk => clk, reset => reset); --
    end block;
    phi_stmt_3026_req_16325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1969), ack => phi_stmt_3026_req_0); -- 
    -- CP-element group 1970 join  transition  bypass 
    -- predecessors 1963 1969 
    -- successors 1981 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_bbx_xnphx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1970: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1970"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1963) & cp_elements(1969);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1970), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1971 fork  transition  bypass 
    -- predecessors 49 
    -- successors 1972 1976 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/$entry
      -- 
    cp_elements(1971) <= cp_elements(49);
    -- CP-element group 1972 fork  transition  bypass 
    -- predecessors 1971 
    -- successors 1973 1974 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/$entry
      -- 
    cp_elements(1972) <= cp_elements(1971);
    -- CP-element group 1973 transition  bypass 
    -- predecessors 1972 
    -- successors 1975 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Sample/ra
      -- 
    cp_elements(1973) <= cp_elements(1972);
    -- CP-element group 1974 transition  bypass 
    -- predecessors 1972 
    -- successors 1975 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/Update/ca
      -- 
    cp_elements(1974) <= cp_elements(1972);
    -- CP-element group 1975 join  transition  output  bypass 
    -- predecessors 1973 1974 
    -- successors 1980 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_sources/type_cast_3022/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3019/phi_stmt_3019_req
      -- 
    cp_element_group_1975: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1975"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1973) & cp_elements(1974);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1975), clk => clk, reset => reset); --
    end block;
    phi_stmt_3019_req_16351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1975), ack => phi_stmt_3019_req_1); -- 
    -- CP-element group 1976 fork  transition  bypass 
    -- predecessors 1971 
    -- successors 1977 1978 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/$entry
      -- 
    cp_elements(1976) <= cp_elements(1971);
    -- CP-element group 1977 transition  bypass 
    -- predecessors 1976 
    -- successors 1979 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Sample/ra
      -- 
    cp_elements(1977) <= cp_elements(1976);
    -- CP-element group 1978 transition  bypass 
    -- predecessors 1976 
    -- successors 1979 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/Update/ca
      -- 
    cp_elements(1978) <= cp_elements(1976);
    -- CP-element group 1979 join  transition  output  bypass 
    -- predecessors 1977 1978 
    -- successors 1980 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_sources/type_cast_3029/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/phi_stmt_3026/phi_stmt_3026_req
      -- 
    cp_element_group_1979: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1979"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1977) & cp_elements(1978);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1979), clk => clk, reset => reset); --
    end block;
    phi_stmt_3026_req_16374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1979), ack => phi_stmt_3026_req_1); -- 
    -- CP-element group 1980 join  transition  bypass 
    -- predecessors 1975 1979 
    -- successors 1981 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xix_xpreheader_bbx_xnphx_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_1980: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1980"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1975) & cp_elements(1979);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1980), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1981 merge  place  bypass 
    -- predecessors 1970 1980 
    -- successors 1982 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3018_PhiReqMerge
      -- 
    cp_elements(1981) <= OrReduce(cp_elements(1970) & cp_elements(1980));
    -- CP-element group 1982 fork  transition  bypass 
    -- predecessors 1981 
    -- successors 1983 1984 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3018_PhiAck/$entry
      -- 
    cp_elements(1982) <= cp_elements(1981);
    -- CP-element group 1983 transition  input  bypass 
    -- predecessors 1982 
    -- successors 1985 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3018_PhiAck/phi_stmt_3019_ack
      -- 
    phi_stmt_3019_ack_16379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3019_ack_0, ack => cp_elements(1983)); -- 
    -- CP-element group 1984 transition  input  bypass 
    -- predecessors 1982 
    -- successors 1985 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3018_PhiAck/phi_stmt_3026_ack
      -- 
    phi_stmt_3026_ack_16380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3026_ack_0, ack => cp_elements(1984)); -- 
    -- CP-element group 1985 join  transition  bypass 
    -- predecessors 1983 1984 
    -- successors 50 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3018_PhiAck/$exit
      -- 
    cp_element_group_1985: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1985"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1983) & cp_elements(1984);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1985), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1986 fork  transition  bypass 
    -- predecessors 908 
    -- successors 1987 1993 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/$entry
      -- 
    cp_elements(1986) <= cp_elements(908);
    -- CP-element group 1987 fork  transition  bypass 
    -- predecessors 1986 
    -- successors 1988 1990 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/$entry
      -- 
    cp_elements(1987) <= cp_elements(1986);
    -- CP-element group 1988 transition  output  bypass 
    -- predecessors 1987 
    -- successors 1989 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Sample/rr
      -- 
    cp_elements(1988) <= cp_elements(1987);
    rr_16403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1988), ack => type_cast_3061_inst_req_0); -- 
    -- CP-element group 1989 transition  input  bypass 
    -- predecessors 1988 
    -- successors 1992 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Sample/ra
      -- 
    ra_16404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3061_inst_ack_0, ack => cp_elements(1989)); -- 
    -- CP-element group 1990 transition  output  bypass 
    -- predecessors 1987 
    -- successors 1991 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Update/cr
      -- 
    cp_elements(1990) <= cp_elements(1987);
    cr_16408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1990), ack => type_cast_3061_inst_req_1); -- 
    -- CP-element group 1991 transition  input  bypass 
    -- predecessors 1990 
    -- successors 1992 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/Update/ca
      -- 
    ca_16409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3061_inst_ack_1, ack => cp_elements(1991)); -- 
    -- CP-element group 1992 join  transition  output  bypass 
    -- predecessors 1989 1991 
    -- successors 1999 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_sources/type_cast_3061/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3058/phi_stmt_3058_req
      -- 
    cp_element_group_1992: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1992"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1989) & cp_elements(1991);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1992), clk => clk, reset => reset); --
    end block;
    phi_stmt_3058_req_16410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1992), ack => phi_stmt_3058_req_0); -- 
    -- CP-element group 1993 fork  transition  bypass 
    -- predecessors 1986 
    -- successors 1994 1996 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/$entry
      -- 
    cp_elements(1993) <= cp_elements(1986);
    -- CP-element group 1994 transition  output  bypass 
    -- predecessors 1993 
    -- successors 1995 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Sample/rr
      -- 
    cp_elements(1994) <= cp_elements(1993);
    rr_16426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1994), ack => type_cast_3065_inst_req_0); -- 
    -- CP-element group 1995 transition  input  bypass 
    -- predecessors 1994 
    -- successors 1998 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Sample/ra
      -- 
    ra_16427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3065_inst_ack_0, ack => cp_elements(1995)); -- 
    -- CP-element group 1996 transition  output  bypass 
    -- predecessors 1993 
    -- successors 1997 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Update/cr
      -- 
    cp_elements(1996) <= cp_elements(1993);
    cr_16431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1996), ack => type_cast_3065_inst_req_1); -- 
    -- CP-element group 1997 transition  input  bypass 
    -- predecessors 1996 
    -- successors 1998 
    -- members (2) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/Update/ca
      -- 
    ca_16432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3065_inst_ack_1, ack => cp_elements(1997)); -- 
    -- CP-element group 1998 join  transition  output  bypass 
    -- predecessors 1995 1997 
    -- successors 1999 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_sources/type_cast_3065/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/phi_stmt_3062/phi_stmt_3062_req
      -- 
    cp_element_group_1998: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1998"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1995) & cp_elements(1997);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1998), clk => clk, reset => reset); --
    end block;
    phi_stmt_3062_req_16433_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1998), ack => phi_stmt_3062_req_0); -- 
    -- CP-element group 1999 join  transition  bypass 
    -- predecessors 1992 1998 
    -- successors 2000 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnphx_xix_xi_xx_x_crit_edgex_xix_xix_xloopexit_PhiReq/$exit
      -- 
    cp_element_group_1999: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_1999"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(1992) & cp_elements(1998);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(1999), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2000 place  bypass 
    -- predecessors 1999 
    -- successors 2001 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3057_PhiReqMerge
      -- 
    cp_elements(2000) <= cp_elements(1999);
    -- CP-element group 2001 fork  transition  bypass 
    -- predecessors 2000 
    -- successors 2002 2003 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3057_PhiAck/$entry
      -- 
    cp_elements(2001) <= cp_elements(2000);
    -- CP-element group 2002 transition  input  bypass 
    -- predecessors 2001 
    -- successors 2004 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3057_PhiAck/phi_stmt_3058_ack
      -- 
    phi_stmt_3058_ack_16438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3058_ack_0, ack => cp_elements(2002)); -- 
    -- CP-element group 2003 transition  input  bypass 
    -- predecessors 2001 
    -- successors 2004 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3057_PhiAck/phi_stmt_3062_ack
      -- 
    phi_stmt_3062_ack_16439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3062_ack_0, ack => cp_elements(2003)); -- 
    -- CP-element group 2004 join  transition  bypass 
    -- predecessors 2002 2003 
    -- successors 52 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3057_PhiAck/$exit
      -- 
    cp_element_group_2004: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2004"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2002) & cp_elements(2003);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2004), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2005 fork  transition  bypass 
    -- predecessors 886 
    -- successors 2006 2010 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2005) <= cp_elements(886);
    -- CP-element group 2006 fork  transition  bypass 
    -- predecessors 2005 
    -- successors 2007 2008 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/$entry
      -- 
    cp_elements(2006) <= cp_elements(2005);
    -- CP-element group 2007 transition  bypass 
    -- predecessors 2006 
    -- successors 2009 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/ra
      -- 
    cp_elements(2007) <= cp_elements(2006);
    -- CP-element group 2008 transition  bypass 
    -- predecessors 2006 
    -- successors 2009 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/ca
      -- 
    cp_elements(2008) <= cp_elements(2006);
    -- CP-element group 2009 join  transition  output  bypass 
    -- predecessors 2007 2008 
    -- successors 2014 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_req
      -- 
    cp_element_group_2009: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2009"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2007) & cp_elements(2008);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2009), clk => clk, reset => reset); --
    end block;
    phi_stmt_3069_req_16465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2009), ack => phi_stmt_3069_req_0); -- 
    -- CP-element group 2010 fork  transition  bypass 
    -- predecessors 2005 
    -- successors 2011 2012 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/$entry
      -- 
    cp_elements(2010) <= cp_elements(2005);
    -- CP-element group 2011 transition  bypass 
    -- predecessors 2010 
    -- successors 2013 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/ra
      -- 
    cp_elements(2011) <= cp_elements(2010);
    -- CP-element group 2012 transition  bypass 
    -- predecessors 2010 
    -- successors 2013 
    -- members (4) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/ca
      -- 
    cp_elements(2012) <= cp_elements(2010);
    -- CP-element group 2013 join  transition  output  bypass 
    -- predecessors 2011 2012 
    -- successors 2014 
    -- members (5) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_req
      -- 
    cp_element_group_2013: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2013"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2011) & cp_elements(2012);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2013), clk => clk, reset => reset); --
    end block;
    phi_stmt_3076_req_16488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2013), ack => phi_stmt_3076_req_0); -- 
    -- CP-element group 2014 join  transition  bypass 
    -- predecessors 2009 2013 
    -- successors 2029 
    -- members (1) 
      -- 	branch_block_stmt_1659/bbx_xnph7x_xix_xi_xx_x_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2014: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2014"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2009) & cp_elements(2013);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2014), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2015 fork  transition  bypass 
    -- predecessors 52 
    -- successors 2016 2022 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/$entry
      -- 
    cp_elements(2015) <= cp_elements(52);
    -- CP-element group 2016 fork  transition  bypass 
    -- predecessors 2015 
    -- successors 2017 2019 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/$entry
      -- 
    cp_elements(2016) <= cp_elements(2015);
    -- CP-element group 2017 transition  output  bypass 
    -- predecessors 2016 
    -- successors 2018 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/rr
      -- 
    cp_elements(2017) <= cp_elements(2016);
    rr_16507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2017), ack => type_cast_3075_inst_req_0); -- 
    -- CP-element group 2018 transition  input  bypass 
    -- predecessors 2017 
    -- successors 2021 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Sample/ra
      -- 
    ra_16508_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3075_inst_ack_0, ack => cp_elements(2018)); -- 
    -- CP-element group 2019 transition  output  bypass 
    -- predecessors 2016 
    -- successors 2020 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/cr
      -- 
    cp_elements(2019) <= cp_elements(2016);
    cr_16512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2019), ack => type_cast_3075_inst_req_1); -- 
    -- CP-element group 2020 transition  input  bypass 
    -- predecessors 2019 
    -- successors 2021 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/Update/ca
      -- 
    ca_16513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3075_inst_ack_1, ack => cp_elements(2020)); -- 
    -- CP-element group 2021 join  transition  output  bypass 
    -- predecessors 2018 2020 
    -- successors 2028 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_sources/type_cast_3075/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3069/phi_stmt_3069_req
      -- 
    cp_element_group_2021: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2021"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2018) & cp_elements(2020);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2021), clk => clk, reset => reset); --
    end block;
    phi_stmt_3069_req_16514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2021), ack => phi_stmt_3069_req_1); -- 
    -- CP-element group 2022 fork  transition  bypass 
    -- predecessors 2015 
    -- successors 2023 2025 
    -- members (4) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/$entry
      -- 
    cp_elements(2022) <= cp_elements(2015);
    -- CP-element group 2023 transition  output  bypass 
    -- predecessors 2022 
    -- successors 2024 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/rr
      -- 
    cp_elements(2023) <= cp_elements(2022);
    rr_16530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2023), ack => type_cast_3082_inst_req_0); -- 
    -- CP-element group 2024 transition  input  bypass 
    -- predecessors 2023 
    -- successors 2027 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Sample/ra
      -- 
    ra_16531_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3082_inst_ack_0, ack => cp_elements(2024)); -- 
    -- CP-element group 2025 transition  output  bypass 
    -- predecessors 2022 
    -- successors 2026 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/cr
      -- 
    cp_elements(2025) <= cp_elements(2022);
    cr_16535_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2025), ack => type_cast_3082_inst_req_1); -- 
    -- CP-element group 2026 transition  input  bypass 
    -- predecessors 2025 
    -- successors 2027 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/Update/ca
      -- 
    ca_16536_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3082_inst_ack_1, ack => cp_elements(2026)); -- 
    -- CP-element group 2027 join  transition  output  bypass 
    -- predecessors 2024 2026 
    -- successors 2028 
    -- members (5) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_sources/type_cast_3082/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/phi_stmt_3076/phi_stmt_3076_req
      -- 
    cp_element_group_2027: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2027"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2024) & cp_elements(2026);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2027), clk => clk, reset => reset); --
    end block;
    phi_stmt_3076_req_16537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2027), ack => phi_stmt_3076_req_1); -- 
    -- CP-element group 2028 join  transition  bypass 
    -- predecessors 2021 2027 
    -- successors 2029 
    -- members (1) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xix_xloopexit_xx_x_crit_edgex_xix_xi_PhiReq/$exit
      -- 
    cp_element_group_2028: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2028"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2021) & cp_elements(2027);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2028), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2029 merge  place  bypass 
    -- predecessors 2014 2028 
    -- successors 2030 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3068_PhiReqMerge
      -- 
    cp_elements(2029) <= OrReduce(cp_elements(2014) & cp_elements(2028));
    -- CP-element group 2030 fork  transition  bypass 
    -- predecessors 2029 
    -- successors 2031 2032 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3068_PhiAck/$entry
      -- 
    cp_elements(2030) <= cp_elements(2029);
    -- CP-element group 2031 transition  input  bypass 
    -- predecessors 2030 
    -- successors 2033 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3068_PhiAck/phi_stmt_3069_ack
      -- 
    phi_stmt_3069_ack_16542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3069_ack_0, ack => cp_elements(2031)); -- 
    -- CP-element group 2032 transition  input  bypass 
    -- predecessors 2030 
    -- successors 2033 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3068_PhiAck/phi_stmt_3076_ack
      -- 
    phi_stmt_3076_ack_16543_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3076_ack_0, ack => cp_elements(2032)); -- 
    -- CP-element group 2033 join  transition  bypass 
    -- predecessors 2031 2032 
    -- successors 53 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3068_PhiAck/$exit
      -- 
    cp_element_group_2033: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2033"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2031) & cp_elements(2032);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2033), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2034 transition  output  bypass 
    -- predecessors 930 
    -- successors 2035 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Sample/rr
      -- 
    cp_elements(2034) <= cp_elements(930);
    rr_16566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2034), ack => type_cast_3110_inst_req_0); -- 
    -- CP-element group 2035 transition  input  bypass 
    -- predecessors 2034 
    -- successors 2038 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Sample/ra
      -- 
    ra_16567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3110_inst_ack_0, ack => cp_elements(2035)); -- 
    -- CP-element group 2036 transition  output  bypass 
    -- predecessors 930 
    -- successors 2037 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Update/cr
      -- 
    cp_elements(2036) <= cp_elements(930);
    cr_16571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2036), ack => type_cast_3110_inst_req_1); -- 
    -- CP-element group 2037 transition  input  bypass 
    -- predecessors 2036 
    -- successors 2038 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/Update/ca
      -- 
    ca_16572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3110_inst_ack_1, ack => cp_elements(2037)); -- 
    -- CP-element group 2038 join  transition  place  output  bypass 
    -- predecessors 2035 2037 
    -- successors 2039 
    -- members (8) 
      -- 	branch_block_stmt_1659/merge_stmt_3106_PhiReqMerge
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_sources/type_cast_3110/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_x_crit_edgex_xix_xi_udiv32x_xexitx_xpreheaderx_xi_PhiReq/phi_stmt_3107/phi_stmt_3107_req
      -- 	branch_block_stmt_1659/merge_stmt_3106_PhiAck/$entry
      -- 
    cp_element_group_2038: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2038"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2035) & cp_elements(2037);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2038), clk => clk, reset => reset); --
    end block;
    phi_stmt_3107_req_16573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2038), ack => phi_stmt_3107_req_0); -- 
    -- CP-element group 2039 transition  input  bypass 
    -- predecessors 2038 
    -- successors 55 
    -- members (2) 
      -- 	branch_block_stmt_1659/merge_stmt_3106_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3106_PhiAck/phi_stmt_3107_ack
      -- 
    phi_stmt_3107_ack_16578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3107_ack_0, ack => cp_elements(2039)); -- 
    -- CP-element group 2040 fork  transition  bypass 
    -- predecessors 1004 
    -- successors 2041 2047 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/$entry
      -- 
    cp_elements(2040) <= cp_elements(1004);
    -- CP-element group 2041 fork  transition  bypass 
    -- predecessors 2040 
    -- successors 2042 2044 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/$entry
      -- 
    cp_elements(2041) <= cp_elements(2040);
    -- CP-element group 2042 transition  output  bypass 
    -- predecessors 2041 
    -- successors 2043 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/rr
      -- 
    cp_elements(2042) <= cp_elements(2041);
    rr_16609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2042), ack => type_cast_3173_inst_req_0); -- 
    -- CP-element group 2043 transition  input  bypass 
    -- predecessors 2042 
    -- successors 2046 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/ra
      -- 
    ra_16610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3173_inst_ack_0, ack => cp_elements(2043)); -- 
    -- CP-element group 2044 transition  output  bypass 
    -- predecessors 2041 
    -- successors 2045 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/cr
      -- 
    cp_elements(2044) <= cp_elements(2041);
    cr_16614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2044), ack => type_cast_3173_inst_req_1); -- 
    -- CP-element group 2045 transition  input  bypass 
    -- predecessors 2044 
    -- successors 2046 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/ca
      -- 
    ca_16615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3173_inst_ack_1, ack => cp_elements(2045)); -- 
    -- CP-element group 2046 join  transition  output  bypass 
    -- predecessors 2043 2045 
    -- successors 2059 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_req
      -- 
    cp_element_group_2046: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2046"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2043) & cp_elements(2045);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2046), clk => clk, reset => reset); --
    end block;
    phi_stmt_3170_req_16616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2046), ack => phi_stmt_3170_req_0); -- 
    -- CP-element group 2047 fork  transition  bypass 
    -- predecessors 2040 
    -- successors 2048 2054 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/$entry
      -- 
    cp_elements(2047) <= cp_elements(2040);
    -- CP-element group 2048 fork  transition  bypass 
    -- predecessors 2047 
    -- successors 2049 2051 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/$entry
      -- 
    cp_elements(2048) <= cp_elements(2047);
    -- CP-element group 2049 transition  output  bypass 
    -- predecessors 2048 
    -- successors 2050 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/rr
      -- 
    cp_elements(2049) <= cp_elements(2048);
    rr_16632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2049), ack => type_cast_3180_inst_req_0); -- 
    -- CP-element group 2050 transition  input  bypass 
    -- predecessors 2049 
    -- successors 2053 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/ra
      -- 
    ra_16633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3180_inst_ack_0, ack => cp_elements(2050)); -- 
    -- CP-element group 2051 transition  output  bypass 
    -- predecessors 2048 
    -- successors 2052 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/cr
      -- 
    cp_elements(2051) <= cp_elements(2048);
    cr_16637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2051), ack => type_cast_3180_inst_req_1); -- 
    -- CP-element group 2052 transition  input  bypass 
    -- predecessors 2051 
    -- successors 2053 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/ca
      -- 
    ca_16638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3180_inst_ack_1, ack => cp_elements(2052)); -- 
    -- CP-element group 2053 join  transition  bypass 
    -- predecessors 2050 2052 
    -- successors 2058 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/$exit
      -- 
    cp_element_group_2053: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2053"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2050) & cp_elements(2052);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2053), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2054 fork  transition  bypass 
    -- predecessors 2047 
    -- successors 2055 2056 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/$entry
      -- 
    cp_elements(2054) <= cp_elements(2047);
    -- CP-element group 2055 transition  bypass 
    -- predecessors 2054 
    -- successors 2057 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/ra
      -- 
    cp_elements(2055) <= cp_elements(2054);
    -- CP-element group 2056 transition  bypass 
    -- predecessors 2054 
    -- successors 2057 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/ca
      -- 
    cp_elements(2056) <= cp_elements(2054);
    -- CP-element group 2057 join  transition  bypass 
    -- predecessors 2055 2056 
    -- successors 2058 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/$exit
      -- 
    cp_element_group_2057: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2057"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2055) & cp_elements(2056);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2057), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2058 join  transition  output  bypass 
    -- predecessors 2053 2057 
    -- successors 2059 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_req
      -- 
    cp_element_group_2058: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2058"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2053) & cp_elements(2057);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2058), clk => clk, reset => reset); --
    end block;
    phi_stmt_3177_req_16655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2058), ack => phi_stmt_3177_req_0); -- 
    -- CP-element group 2059 join  transition  bypass 
    -- predecessors 2046 2058 
    -- successors 2078 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xi_PhiReq/$exit
      -- 
    cp_element_group_2059: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2059"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2046) & cp_elements(2058);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2059), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2060 fork  transition  bypass 
    -- predecessors 57 
    -- successors 2061 2065 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/$entry
      -- 
    cp_elements(2060) <= cp_elements(57);
    -- CP-element group 2061 fork  transition  bypass 
    -- predecessors 2060 
    -- successors 2062 2063 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/$entry
      -- 
    cp_elements(2061) <= cp_elements(2060);
    -- CP-element group 2062 transition  bypass 
    -- predecessors 2061 
    -- successors 2064 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Sample/ra
      -- 
    cp_elements(2062) <= cp_elements(2061);
    -- CP-element group 2063 transition  bypass 
    -- predecessors 2061 
    -- successors 2064 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/Update/ca
      -- 
    cp_elements(2063) <= cp_elements(2061);
    -- CP-element group 2064 join  transition  output  bypass 
    -- predecessors 2062 2063 
    -- successors 2077 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_sources/type_cast_3173/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3170/phi_stmt_3170_req
      -- 
    cp_element_group_2064: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2064"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2062) & cp_elements(2063);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2064), clk => clk, reset => reset); --
    end block;
    phi_stmt_3170_req_16681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2064), ack => phi_stmt_3170_req_1); -- 
    -- CP-element group 2065 fork  transition  bypass 
    -- predecessors 2060 
    -- successors 2066 2070 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/$entry
      -- 
    cp_elements(2065) <= cp_elements(2060);
    -- CP-element group 2066 fork  transition  bypass 
    -- predecessors 2065 
    -- successors 2067 2068 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/$entry
      -- 
    cp_elements(2066) <= cp_elements(2065);
    -- CP-element group 2067 transition  bypass 
    -- predecessors 2066 
    -- successors 2069 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Sample/ra
      -- 
    cp_elements(2067) <= cp_elements(2066);
    -- CP-element group 2068 transition  bypass 
    -- predecessors 2066 
    -- successors 2069 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/Update/ca
      -- 
    cp_elements(2068) <= cp_elements(2066);
    -- CP-element group 2069 join  transition  bypass 
    -- predecessors 2067 2068 
    -- successors 2076 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3180/SplitProtocol/$exit
      -- 
    cp_element_group_2069: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2069"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2067) & cp_elements(2068);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2069), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2070 fork  transition  bypass 
    -- predecessors 2065 
    -- successors 2071 2073 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/$entry
      -- 
    cp_elements(2070) <= cp_elements(2065);
    -- CP-element group 2071 transition  output  bypass 
    -- predecessors 2070 
    -- successors 2072 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/rr
      -- 
    cp_elements(2071) <= cp_elements(2070);
    rr_16713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2071), ack => type_cast_3182_inst_req_0); -- 
    -- CP-element group 2072 transition  input  bypass 
    -- predecessors 2071 
    -- successors 2075 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Sample/ra
      -- 
    ra_16714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3182_inst_ack_0, ack => cp_elements(2072)); -- 
    -- CP-element group 2073 transition  output  bypass 
    -- predecessors 2070 
    -- successors 2074 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/cr
      -- 
    cp_elements(2073) <= cp_elements(2070);
    cr_16718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2073), ack => type_cast_3182_inst_req_1); -- 
    -- CP-element group 2074 transition  input  bypass 
    -- predecessors 2073 
    -- successors 2075 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/Update/ca
      -- 
    ca_16719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3182_inst_ack_1, ack => cp_elements(2074)); -- 
    -- CP-element group 2075 join  transition  bypass 
    -- predecessors 2072 2074 
    -- successors 2076 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/type_cast_3182/SplitProtocol/$exit
      -- 
    cp_element_group_2075: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2075"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2072) & cp_elements(2074);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2075), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2076 join  transition  output  bypass 
    -- predecessors 2069 2075 
    -- successors 2077 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/phi_stmt_3177/phi_stmt_3177_req
      -- 
    cp_element_group_2076: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2076"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2069) & cp_elements(2075);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2076), clk => clk, reset => reset); --
    end block;
    phi_stmt_3177_req_16720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2076), ack => phi_stmt_3177_req_1); -- 
    -- CP-element group 2077 join  transition  bypass 
    -- predecessors 2064 2076 
    -- successors 2078 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xix_xpreheader_udiv32x_xexitx_xi_PhiReq/$exit
      -- 
    cp_element_group_2077: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2077"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2064) & cp_elements(2076);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2077), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2078 merge  place  bypass 
    -- predecessors 2059 2077 
    -- successors 2079 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3169_PhiReqMerge
      -- 
    cp_elements(2078) <= OrReduce(cp_elements(2059) & cp_elements(2077));
    -- CP-element group 2079 fork  transition  bypass 
    -- predecessors 2078 
    -- successors 2080 2081 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3169_PhiAck/$entry
      -- 
    cp_elements(2079) <= cp_elements(2078);
    -- CP-element group 2080 transition  input  bypass 
    -- predecessors 2079 
    -- successors 2082 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3169_PhiAck/phi_stmt_3170_ack
      -- 
    phi_stmt_3170_ack_16725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3170_ack_0, ack => cp_elements(2080)); -- 
    -- CP-element group 2081 transition  input  bypass 
    -- predecessors 2079 
    -- successors 2082 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3169_PhiAck/phi_stmt_3177_ack
      -- 
    phi_stmt_3177_ack_16726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3177_ack_0, ack => cp_elements(2081)); -- 
    -- CP-element group 2082 join  transition  bypass 
    -- predecessors 2080 2081 
    -- successors 58 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3169_PhiAck/$exit
      -- 
    cp_element_group_2082: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2082"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2080) & cp_elements(2081);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2082), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2083 fork  transition  bypass 
    -- predecessors 1006 
    -- successors 2084 2090 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/$entry
      -- 
    cp_elements(2083) <= cp_elements(1006);
    -- CP-element group 2084 fork  transition  bypass 
    -- predecessors 2083 
    -- successors 2085 2087 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/$entry
      -- 
    cp_elements(2084) <= cp_elements(2083);
    -- CP-element group 2085 transition  output  bypass 
    -- predecessors 2084 
    -- successors 2086 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Sample/rr
      -- 
    cp_elements(2085) <= cp_elements(2084);
    rr_16749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2085), ack => type_cast_3235_inst_req_0); -- 
    -- CP-element group 2086 transition  input  bypass 
    -- predecessors 2085 
    -- successors 2089 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Sample/ra
      -- 
    ra_16750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3235_inst_ack_0, ack => cp_elements(2086)); -- 
    -- CP-element group 2087 transition  output  bypass 
    -- predecessors 2084 
    -- successors 2088 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Update/cr
      -- 
    cp_elements(2087) <= cp_elements(2084);
    cr_16754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2087), ack => type_cast_3235_inst_req_1); -- 
    -- CP-element group 2088 transition  input  bypass 
    -- predecessors 2087 
    -- successors 2089 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/Update/ca
      -- 
    ca_16755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3235_inst_ack_1, ack => cp_elements(2088)); -- 
    -- CP-element group 2089 join  transition  output  bypass 
    -- predecessors 2086 2088 
    -- successors 2096 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_sources/type_cast_3235/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3232/phi_stmt_3232_req
      -- 
    cp_element_group_2089: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2089"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2086) & cp_elements(2088);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2089), clk => clk, reset => reset); --
    end block;
    phi_stmt_3232_req_16756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2089), ack => phi_stmt_3232_req_0); -- 
    -- CP-element group 2090 fork  transition  bypass 
    -- predecessors 2083 
    -- successors 2091 2093 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/$entry
      -- 
    cp_elements(2090) <= cp_elements(2083);
    -- CP-element group 2091 transition  output  bypass 
    -- predecessors 2090 
    -- successors 2092 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Sample/rr
      -- 
    cp_elements(2091) <= cp_elements(2090);
    rr_16772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2091), ack => type_cast_3231_inst_req_0); -- 
    -- CP-element group 2092 transition  input  bypass 
    -- predecessors 2091 
    -- successors 2095 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Sample/ra
      -- 
    ra_16773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3231_inst_ack_0, ack => cp_elements(2092)); -- 
    -- CP-element group 2093 transition  output  bypass 
    -- predecessors 2090 
    -- successors 2094 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Update/cr
      -- 
    cp_elements(2093) <= cp_elements(2090);
    cr_16777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2093), ack => type_cast_3231_inst_req_1); -- 
    -- CP-element group 2094 transition  input  bypass 
    -- predecessors 2093 
    -- successors 2095 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/Update/ca
      -- 
    ca_16778_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3231_inst_ack_1, ack => cp_elements(2094)); -- 
    -- CP-element group 2095 join  transition  output  bypass 
    -- predecessors 2092 2094 
    -- successors 2096 
    -- members (5) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_sources/type_cast_3231/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/phi_stmt_3228/phi_stmt_3228_req
      -- 
    cp_element_group_2095: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2095"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2092) & cp_elements(2094);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2095), clk => clk, reset => reset); --
    end block;
    phi_stmt_3228_req_16779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2095), ack => phi_stmt_3228_req_0); -- 
    -- CP-element group 2096 join  transition  bypass 
    -- predecessors 2089 2095 
    -- successors 2097 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xi_udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2096: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2096"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2089) & cp_elements(2095);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2096), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2097 place  bypass 
    -- predecessors 2096 
    -- successors 2098 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3227_PhiReqMerge
      -- 
    cp_elements(2097) <= cp_elements(2096);
    -- CP-element group 2098 fork  transition  bypass 
    -- predecessors 2097 
    -- successors 2099 2100 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3227_PhiAck/$entry
      -- 
    cp_elements(2098) <= cp_elements(2097);
    -- CP-element group 2099 transition  input  bypass 
    -- predecessors 2098 
    -- successors 2101 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3227_PhiAck/phi_stmt_3228_ack
      -- 
    phi_stmt_3228_ack_16784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3228_ack_0, ack => cp_elements(2099)); -- 
    -- CP-element group 2100 transition  input  bypass 
    -- predecessors 2098 
    -- successors 2101 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3227_PhiAck/phi_stmt_3232_ack
      -- 
    phi_stmt_3232_ack_16785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3232_ack_0, ack => cp_elements(2100)); -- 
    -- CP-element group 2101 join  transition  bypass 
    -- predecessors 2099 2100 
    -- successors 60 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3227_PhiAck/$exit
      -- 
    cp_element_group_2101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2099) & cp_elements(2100);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2102 fork  transition  bypass 
    -- predecessors 972 
    -- successors 2103 2115 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/$entry
      -- 
    cp_elements(2102) <= cp_elements(972);
    -- CP-element group 2103 fork  transition  bypass 
    -- predecessors 2102 
    -- successors 2104 2108 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/$entry
      -- 
    cp_elements(2103) <= cp_elements(2102);
    -- CP-element group 2104 fork  transition  bypass 
    -- predecessors 2103 
    -- successors 2105 2106 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/$entry
      -- 
    cp_elements(2104) <= cp_elements(2103);
    -- CP-element group 2105 transition  bypass 
    -- predecessors 2104 
    -- successors 2107 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/ra
      -- 
    cp_elements(2105) <= cp_elements(2104);
    -- CP-element group 2106 transition  bypass 
    -- predecessors 2104 
    -- successors 2107 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/ca
      -- 
    cp_elements(2106) <= cp_elements(2104);
    -- CP-element group 2107 join  transition  bypass 
    -- predecessors 2105 2106 
    -- successors 2114 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/$exit
      -- 
    cp_element_group_2107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2105) & cp_elements(2106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2108 fork  transition  bypass 
    -- predecessors 2103 
    -- successors 2109 2111 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/$entry
      -- 
    cp_elements(2108) <= cp_elements(2103);
    -- CP-element group 2109 transition  output  bypass 
    -- predecessors 2108 
    -- successors 2110 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/rr
      -- 
    cp_elements(2109) <= cp_elements(2108);
    rr_16820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2109), ack => type_cast_3255_inst_req_0); -- 
    -- CP-element group 2110 transition  input  bypass 
    -- predecessors 2109 
    -- successors 2113 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/ra
      -- 
    ra_16821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3255_inst_ack_0, ack => cp_elements(2110)); -- 
    -- CP-element group 2111 transition  output  bypass 
    -- predecessors 2108 
    -- successors 2112 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/cr
      -- 
    cp_elements(2111) <= cp_elements(2108);
    cr_16825_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2111), ack => type_cast_3255_inst_req_1); -- 
    -- CP-element group 2112 transition  input  bypass 
    -- predecessors 2111 
    -- successors 2113 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/ca
      -- 
    ca_16826_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3255_inst_ack_1, ack => cp_elements(2112)); -- 
    -- CP-element group 2113 join  transition  bypass 
    -- predecessors 2110 2112 
    -- successors 2114 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/$exit
      -- 
    cp_element_group_2113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2110) & cp_elements(2112);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2114 join  transition  output  bypass 
    -- predecessors 2107 2113 
    -- successors 2127 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_req
      -- 
    cp_element_group_2114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2107) & cp_elements(2113);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2114), clk => clk, reset => reset); --
    end block;
    phi_stmt_3250_req_16827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2114), ack => phi_stmt_3250_req_1); -- 
    -- CP-element group 2115 fork  transition  bypass 
    -- predecessors 2102 
    -- successors 2116 2120 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/$entry
      -- 
    cp_elements(2115) <= cp_elements(2102);
    -- CP-element group 2116 fork  transition  bypass 
    -- predecessors 2115 
    -- successors 2117 2118 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/$entry
      -- 
    cp_elements(2116) <= cp_elements(2115);
    -- CP-element group 2117 transition  bypass 
    -- predecessors 2116 
    -- successors 2119 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/ra
      -- 
    cp_elements(2117) <= cp_elements(2116);
    -- CP-element group 2118 transition  bypass 
    -- predecessors 2116 
    -- successors 2119 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/ca
      -- 
    cp_elements(2118) <= cp_elements(2116);
    -- CP-element group 2119 join  transition  bypass 
    -- predecessors 2117 2118 
    -- successors 2126 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/$exit
      -- 
    cp_element_group_2119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2117) & cp_elements(2118);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2120 fork  transition  bypass 
    -- predecessors 2115 
    -- successors 2121 2123 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/$entry
      -- 
    cp_elements(2120) <= cp_elements(2115);
    -- CP-element group 2121 transition  output  bypass 
    -- predecessors 2120 
    -- successors 2122 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/rr
      -- 
    cp_elements(2121) <= cp_elements(2120);
    rr_16859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2121), ack => type_cast_3261_inst_req_0); -- 
    -- CP-element group 2122 transition  input  bypass 
    -- predecessors 2121 
    -- successors 2125 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/ra
      -- 
    ra_16860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3261_inst_ack_0, ack => cp_elements(2122)); -- 
    -- CP-element group 2123 transition  output  bypass 
    -- predecessors 2120 
    -- successors 2124 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/cr
      -- 
    cp_elements(2123) <= cp_elements(2120);
    cr_16864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2123), ack => type_cast_3261_inst_req_1); -- 
    -- CP-element group 2124 transition  input  bypass 
    -- predecessors 2123 
    -- successors 2125 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/ca
      -- 
    ca_16865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3261_inst_ack_1, ack => cp_elements(2124)); -- 
    -- CP-element group 2125 join  transition  bypass 
    -- predecessors 2122 2124 
    -- successors 2126 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/$exit
      -- 
    cp_element_group_2125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2122) & cp_elements(2124);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2126 join  transition  output  bypass 
    -- predecessors 2119 2125 
    -- successors 2127 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_req
      -- 
    cp_element_group_2126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2119) & cp_elements(2125);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2126), clk => clk, reset => reset); --
    end block;
    phi_stmt_3256_req_16866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2126), ack => phi_stmt_3256_req_1); -- 
    -- CP-element group 2127 join  transition  bypass 
    -- predecessors 2114 2126 
    -- successors 2154 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xpreheaderx_xi_xx_xcritedgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2114) & cp_elements(2126);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2128 fork  transition  bypass 
    -- predecessors 1016 
    -- successors 2129 2141 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/$entry
      -- 
    cp_elements(2128) <= cp_elements(1016);
    -- CP-element group 2129 fork  transition  bypass 
    -- predecessors 2128 
    -- successors 2130 2136 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/$entry
      -- 
    cp_elements(2129) <= cp_elements(2128);
    -- CP-element group 2130 fork  transition  bypass 
    -- predecessors 2129 
    -- successors 2131 2133 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/$entry
      -- 
    cp_elements(2130) <= cp_elements(2129);
    -- CP-element group 2131 transition  output  bypass 
    -- predecessors 2130 
    -- successors 2132 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/rr
      -- 
    cp_elements(2131) <= cp_elements(2130);
    rr_16885_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2131), ack => type_cast_3253_inst_req_0); -- 
    -- CP-element group 2132 transition  input  bypass 
    -- predecessors 2131 
    -- successors 2135 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Sample/ra
      -- 
    ra_16886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3253_inst_ack_0, ack => cp_elements(2132)); -- 
    -- CP-element group 2133 transition  output  bypass 
    -- predecessors 2130 
    -- successors 2134 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/cr
      -- 
    cp_elements(2133) <= cp_elements(2130);
    cr_16890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2133), ack => type_cast_3253_inst_req_1); -- 
    -- CP-element group 2134 transition  input  bypass 
    -- predecessors 2133 
    -- successors 2135 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/Update/ca
      -- 
    ca_16891_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3253_inst_ack_1, ack => cp_elements(2134)); -- 
    -- CP-element group 2135 join  transition  bypass 
    -- predecessors 2132 2134 
    -- successors 2140 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3253/SplitProtocol/$exit
      -- 
    cp_element_group_2135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2132) & cp_elements(2134);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2136 fork  transition  bypass 
    -- predecessors 2129 
    -- successors 2137 2138 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/$entry
      -- 
    cp_elements(2136) <= cp_elements(2129);
    -- CP-element group 2137 transition  bypass 
    -- predecessors 2136 
    -- successors 2139 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Sample/ra
      -- 
    cp_elements(2137) <= cp_elements(2136);
    -- CP-element group 2138 transition  bypass 
    -- predecessors 2136 
    -- successors 2139 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/Update/ca
      -- 
    cp_elements(2138) <= cp_elements(2136);
    -- CP-element group 2139 join  transition  bypass 
    -- predecessors 2137 2138 
    -- successors 2140 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/type_cast_3255/SplitProtocol/$exit
      -- 
    cp_element_group_2139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2137) & cp_elements(2138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2140 join  transition  output  bypass 
    -- predecessors 2135 2139 
    -- successors 2153 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3250/phi_stmt_3250_req
      -- 
    cp_element_group_2140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2135) & cp_elements(2139);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2140), clk => clk, reset => reset); --
    end block;
    phi_stmt_3250_req_16908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2140), ack => phi_stmt_3250_req_0); -- 
    -- CP-element group 2141 fork  transition  bypass 
    -- predecessors 2128 
    -- successors 2142 2148 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/$entry
      -- 
    cp_elements(2141) <= cp_elements(2128);
    -- CP-element group 2142 fork  transition  bypass 
    -- predecessors 2141 
    -- successors 2143 2145 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/$entry
      -- 
    cp_elements(2142) <= cp_elements(2141);
    -- CP-element group 2143 transition  output  bypass 
    -- predecessors 2142 
    -- successors 2144 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/rr
      -- 
    cp_elements(2143) <= cp_elements(2142);
    rr_16924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2143), ack => type_cast_3259_inst_req_0); -- 
    -- CP-element group 2144 transition  input  bypass 
    -- predecessors 2143 
    -- successors 2147 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Sample/ra
      -- 
    ra_16925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3259_inst_ack_0, ack => cp_elements(2144)); -- 
    -- CP-element group 2145 transition  output  bypass 
    -- predecessors 2142 
    -- successors 2146 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/cr
      -- 
    cp_elements(2145) <= cp_elements(2142);
    cr_16929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2145), ack => type_cast_3259_inst_req_1); -- 
    -- CP-element group 2146 transition  input  bypass 
    -- predecessors 2145 
    -- successors 2147 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/Update/ca
      -- 
    ca_16930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3259_inst_ack_1, ack => cp_elements(2146)); -- 
    -- CP-element group 2147 join  transition  bypass 
    -- predecessors 2144 2146 
    -- successors 2152 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3259/SplitProtocol/$exit
      -- 
    cp_element_group_2147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2144) & cp_elements(2146);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2148 fork  transition  bypass 
    -- predecessors 2141 
    -- successors 2149 2150 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/$entry
      -- 
    cp_elements(2148) <= cp_elements(2141);
    -- CP-element group 2149 transition  bypass 
    -- predecessors 2148 
    -- successors 2151 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Sample/ra
      -- 
    cp_elements(2149) <= cp_elements(2148);
    -- CP-element group 2150 transition  bypass 
    -- predecessors 2148 
    -- successors 2151 
    -- members (4) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/Update/ca
      -- 
    cp_elements(2150) <= cp_elements(2148);
    -- CP-element group 2151 join  transition  bypass 
    -- predecessors 2149 2150 
    -- successors 2152 
    -- members (2) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/type_cast_3261/SplitProtocol/$exit
      -- 
    cp_element_group_2151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2149) & cp_elements(2150);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2152 join  transition  output  bypass 
    -- predecessors 2147 2151 
    -- successors 2153 
    -- members (3) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_sources/$exit
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/phi_stmt_3256/phi_stmt_3256_req
      -- 
    cp_element_group_2152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2147) & cp_elements(2151);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2152), clk => clk, reset => reset); --
    end block;
    phi_stmt_3256_req_16947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2152), ack => phi_stmt_3256_req_0); -- 
    -- CP-element group 2153 join  transition  bypass 
    -- predecessors 2140 2152 
    -- successors 2154 
    -- members (1) 
      -- 	branch_block_stmt_1659/udiv32x_xexitx_xx_xcritedge_crit_edgex_xi_xx_xcritedgex_xi_PhiReq/$exit
      -- 
    cp_element_group_2153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2140) & cp_elements(2152);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2154 merge  place  bypass 
    -- predecessors 2127 2153 
    -- successors 2155 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3249_PhiReqMerge
      -- 
    cp_elements(2154) <= OrReduce(cp_elements(2127) & cp_elements(2153));
    -- CP-element group 2155 fork  transition  bypass 
    -- predecessors 2154 
    -- successors 2156 2157 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3249_PhiAck/$entry
      -- 
    cp_elements(2155) <= cp_elements(2154);
    -- CP-element group 2156 transition  input  bypass 
    -- predecessors 2155 
    -- successors 2158 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3249_PhiAck/phi_stmt_3250_ack
      -- 
    phi_stmt_3250_ack_16952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3250_ack_0, ack => cp_elements(2156)); -- 
    -- CP-element group 2157 transition  input  bypass 
    -- predecessors 2155 
    -- successors 2158 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3249_PhiAck/phi_stmt_3256_ack
      -- 
    phi_stmt_3256_ack_16953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3256_ack_0, ack => cp_elements(2157)); -- 
    -- CP-element group 2158 join  transition  bypass 
    -- predecessors 2156 2157 
    -- successors 61 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3249_PhiAck/$exit
      -- 
    cp_element_group_2158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2156) & cp_elements(2157);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2159 transition  bypass 
    -- predecessors 855 
    -- successors 2161 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/rr
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/ra
      -- 
    cp_elements(2159) <= cp_elements(855);
    -- CP-element group 2160 transition  bypass 
    -- predecessors 855 
    -- successors 2161 
    -- members (4) 
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/cr
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/ca
      -- 
    cp_elements(2160) <= cp_elements(855);
    -- CP-element group 2161 join  transition  output  bypass 
    -- predecessors 2159 2160 
    -- successors 2167 
    -- members (6) 
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/bb_46_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_req
      -- 
    cp_element_group_2161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2159) & cp_elements(2160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2161), clk => clk, reset => reset); --
    end block;
    phi_stmt_3297_req_16979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2161), ack => phi_stmt_3297_req_1); -- 
    -- CP-element group 2162 transition  output  bypass 
    -- predecessors 1040 
    -- successors 2163 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/rr
      -- 
    cp_elements(2162) <= cp_elements(1040);
    rr_16998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2162), ack => type_cast_3300_inst_req_0); -- 
    -- CP-element group 2163 transition  input  bypass 
    -- predecessors 2162 
    -- successors 2166 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Sample/ra
      -- 
    ra_16999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3300_inst_ack_0, ack => cp_elements(2163)); -- 
    -- CP-element group 2164 transition  output  bypass 
    -- predecessors 1040 
    -- successors 2165 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/$entry
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/cr
      -- 
    cp_elements(2164) <= cp_elements(1040);
    cr_17003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2164), ack => type_cast_3300_inst_req_1); -- 
    -- CP-element group 2165 transition  input  bypass 
    -- predecessors 2164 
    -- successors 2166 
    -- members (2) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/Update/ca
      -- 
    ca_17004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3300_inst_ack_1, ack => cp_elements(2165)); -- 
    -- CP-element group 2166 join  transition  output  bypass 
    -- predecessors 2163 2165 
    -- successors 2167 
    -- members (6) 
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_sources/type_cast_3300/SplitProtocol/$exit
      -- 	branch_block_stmt_1659/xx_xcritedgex_xi_fdiv32x_xexit_PhiReq/phi_stmt_3297/phi_stmt_3297_req
      -- 
    cp_element_group_2166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 21) := "cp_element_group_2166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cp_elements(2163) & cp_elements(2165);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cp_elements(2166), clk => clk, reset => reset); --
    end block;
    phi_stmt_3297_req_17005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2166), ack => phi_stmt_3297_req_0); -- 
    -- CP-element group 2167 merge  place  bypass 
    -- predecessors 2161 2166 
    -- successors 2168 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3296_PhiReqMerge
      -- 
    cp_elements(2167) <= OrReduce(cp_elements(2161) & cp_elements(2166));
    -- CP-element group 2168 transition  bypass 
    -- predecessors 2167 
    -- successors 2169 
    -- members (1) 
      -- 	branch_block_stmt_1659/merge_stmt_3296_PhiAck/$entry
      -- 
    cp_elements(2168) <= cp_elements(2167);
    -- CP-element group 2169 transition  place  input  bypass 
    -- predecessors 2168 
    -- successors 1041 
    -- members (4) 
      -- 	branch_block_stmt_1659/assign_stmt_3307__entry__
      -- 	branch_block_stmt_1659/merge_stmt_3296__exit__
      -- 	branch_block_stmt_1659/merge_stmt_3296_PhiAck/$exit
      -- 	branch_block_stmt_1659/merge_stmt_3296_PhiAck/phi_stmt_3297_ack
      -- 
    phi_stmt_3297_ack_17010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3297_ack_0, ack => cp_elements(2169)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal curr_quotientx_x02x_xix_xi_3026 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x02x_xix_xix_xi7_2098 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x02x_xix_xix_xi_2543 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xi_3076 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xix_xi10_2147 : std_logic_vector(31 downto 0);
    signal curr_quotientx_x0x_xlcssax_xix_xix_xi_2592 : std_logic_vector(31 downto 0);
    signal expr_2047_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2047_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_2050_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2050_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_2492_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2492_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_2495_wire_constant : std_logic_vector(31 downto 0);
    signal expr_2495_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expx_x0x_xlcssax_xi_3250 : std_logic_vector(31 downto 0);
    signal expx_x0x_xlcssax_xix_xi26_2326 : std_logic_vector(31 downto 0);
    signal expx_x0x_xlcssax_xix_xi_2771 : std_logic_vector(31 downto 0);
    signal flux_rotor_lpf_prevx_x0_1662 : std_logic_vector(31 downto 0);
    signal flux_rotor_prevx_x0_1690 : std_logic_vector(31 downto 0);
    signal iNsTr_100_2878 : std_logic_vector(0 downto 0);
    signal iNsTr_104_2651 : std_logic_vector(31 downto 0);
    signal iNsTr_105_2657 : std_logic_vector(0 downto 0);
    signal iNsTr_106_2665 : std_logic_vector(0 downto 0);
    signal iNsTr_108_2077 : std_logic_vector(31 downto 0);
    signal iNsTr_109_2082 : std_logic_vector(0 downto 0);
    signal iNsTr_10_1733 : std_logic_vector(31 downto 0);
    signal iNsTr_112_2344 : std_logic_vector(31 downto 0);
    signal iNsTr_113_2350 : std_logic_vector(31 downto 0);
    signal iNsTr_114_2356 : std_logic_vector(31 downto 0);
    signal iNsTr_115_2361 : std_logic_vector(31 downto 0);
    signal iNsTr_116_2366 : std_logic_vector(31 downto 0);
    signal iNsTr_118_2969 : std_logic_vector(31 downto 0);
    signal iNsTr_119_2975 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1738 : std_logic_vector(0 downto 0);
    signal iNsTr_120_2981 : std_logic_vector(31 downto 0);
    signal iNsTr_122_2928 : std_logic_vector(0 downto 0);
    signal iNsTr_125_2522 : std_logic_vector(31 downto 0);
    signal iNsTr_126_2527 : std_logic_vector(0 downto 0);
    signal iNsTr_129_2789 : std_logic_vector(31 downto 0);
    signal iNsTr_130_2795 : std_logic_vector(31 downto 0);
    signal iNsTr_131_2801 : std_logic_vector(31 downto 0);
    signal iNsTr_132_2806 : std_logic_vector(31 downto 0);
    signal iNsTr_133_2811 : std_logic_vector(31 downto 0);
    signal iNsTr_136_2159 : std_logic_vector(31 downto 0);
    signal iNsTr_137_2164 : std_logic_vector(31 downto 0);
    signal iNsTr_138_2169 : std_logic_vector(0 downto 0);
    signal iNsTr_13_1750 : std_logic_vector(63 downto 0);
    signal iNsTr_140_2235 : std_logic_vector(31 downto 0);
    signal iNsTr_141_2254 : std_logic_vector(31 downto 0);
    signal iNsTr_142_2260 : std_logic_vector(31 downto 0);
    signal iNsTr_143_2266 : std_logic_vector(0 downto 0);
    signal iNsTr_144_2274 : std_logic_vector(0 downto 0);
    signal iNsTr_146_3003 : std_logic_vector(31 downto 0);
    signal iNsTr_147_3009 : std_logic_vector(0 downto 0);
    signal iNsTr_149_2941 : std_logic_vector(0 downto 0);
    signal iNsTr_14_1756 : std_logic_vector(63 downto 0);
    signal iNsTr_152_2604 : std_logic_vector(31 downto 0);
    signal iNsTr_153_2609 : std_logic_vector(31 downto 0);
    signal iNsTr_154_2614 : std_logic_vector(0 downto 0);
    signal iNsTr_156_2680 : std_logic_vector(31 downto 0);
    signal iNsTr_157_2699 : std_logic_vector(31 downto 0);
    signal iNsTr_158_2705 : std_logic_vector(31 downto 0);
    signal iNsTr_159_2711 : std_logic_vector(0 downto 0);
    signal iNsTr_15_1760 : std_logic_vector(31 downto 0);
    signal iNsTr_160_2719 : std_logic_vector(0 downto 0);
    signal iNsTr_162_2111 : std_logic_vector(31 downto 0);
    signal iNsTr_163_2117 : std_logic_vector(31 downto 0);
    signal iNsTr_164_2122 : std_logic_vector(0 downto 0);
    signal iNsTr_169_3088 : std_logic_vector(31 downto 0);
    signal iNsTr_170_3093 : std_logic_vector(31 downto 0);
    signal iNsTr_171_3099 : std_logic_vector(0 downto 0);
    signal iNsTr_173_3297 : std_logic_vector(31 downto 0);
    signal iNsTr_17_1767 : std_logic_vector(0 downto 0);
    signal iNsTr_183_2556 : std_logic_vector(31 downto 0);
    signal iNsTr_184_2562 : std_logic_vector(31 downto 0);
    signal iNsTr_185_2567 : std_logic_vector(0 downto 0);
    signal iNsTr_190_3039 : std_logic_vector(31 downto 0);
    signal iNsTr_191_3045 : std_logic_vector(31 downto 0);
    signal iNsTr_192_3050 : std_logic_vector(0 downto 0);
    signal iNsTr_194_3117 : std_logic_vector(31 downto 0);
    signal iNsTr_195_3123 : std_logic_vector(31 downto 0);
    signal iNsTr_196_3129 : std_logic_vector(31 downto 0);
    signal iNsTr_197_3135 : std_logic_vector(31 downto 0);
    signal iNsTr_198_3141 : std_logic_vector(31 downto 0);
    signal iNsTr_199_3147 : std_logic_vector(0 downto 0);
    signal iNsTr_19_1805 : std_logic_vector(31 downto 0);
    signal iNsTr_200_3155 : std_logic_vector(0 downto 0);
    signal iNsTr_205_3268 : std_logic_vector(31 downto 0);
    signal iNsTr_206_3274 : std_logic_vector(31 downto 0);
    signal iNsTr_207_3280 : std_logic_vector(31 downto 0);
    signal iNsTr_208_3285 : std_logic_vector(31 downto 0);
    signal iNsTr_209_3290 : std_logic_vector(31 downto 0);
    signal iNsTr_20_1810 : std_logic_vector(31 downto 0);
    signal iNsTr_211_3170 : std_logic_vector(31 downto 0);
    signal iNsTr_212_3189 : std_logic_vector(31 downto 0);
    signal iNsTr_213_3195 : std_logic_vector(31 downto 0);
    signal iNsTr_214_3201 : std_logic_vector(0 downto 0);
    signal iNsTr_215_3209 : std_logic_vector(0 downto 0);
    signal iNsTr_21_1815 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1820 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1826 : std_logic_vector(31 downto 0);
    signal iNsTr_24_1831 : std_logic_vector(31 downto 0);
    signal iNsTr_25_1835 : std_logic_vector(63 downto 0);
    signal iNsTr_26_1841 : std_logic_vector(0 downto 0);
    signal iNsTr_28_1778 : std_logic_vector(63 downto 0);
    signal iNsTr_29_1784 : std_logic_vector(63 downto 0);
    signal iNsTr_2_1721 : std_logic_vector(31 downto 0);
    signal iNsTr_30_1788 : std_logic_vector(31 downto 0);
    signal iNsTr_32_1880 : std_logic_vector(31 downto 0);
    signal iNsTr_33_1885 : std_logic_vector(31 downto 0);
    signal iNsTr_34_1891 : std_logic_vector(0 downto 0);
    signal iNsTr_36_1854 : std_logic_vector(0 downto 0);
    signal iNsTr_38_1936 : std_logic_vector(31 downto 0);
    signal iNsTr_39_1941 : std_logic_vector(31 downto 0);
    signal iNsTr_40_1947 : std_logic_vector(31 downto 0);
    signal iNsTr_41_1961 : std_logic_vector(0 downto 0);
    signal iNsTr_43_1904 : std_logic_vector(0 downto 0);
    signal iNsTr_46_2373 : std_logic_vector(31 downto 0);
    signal iNsTr_47_2385 : std_logic_vector(31 downto 0);
    signal iNsTr_48_2391 : std_logic_vector(31 downto 0);
    signal iNsTr_49_2396 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1724 : std_logic_vector(31 downto 0);
    signal iNsTr_50_2406 : std_logic_vector(0 downto 0);
    signal iNsTr_52_1974 : std_logic_vector(31 downto 0);
    signal iNsTr_53_1980 : std_logic_vector(31 downto 0);
    signal iNsTr_54_1986 : std_logic_vector(31 downto 0);
    signal iNsTr_55_1992 : std_logic_vector(31 downto 0);
    signal iNsTr_56_1998 : std_logic_vector(31 downto 0);
    signal iNsTr_57_2004 : std_logic_vector(31 downto 0);
    signal iNsTr_58_2010 : std_logic_vector(31 downto 0);
    signal iNsTr_59_2016 : std_logic_vector(31 downto 0);
    signal iNsTr_60_2022 : std_logic_vector(31 downto 0);
    signal iNsTr_61_2028 : std_logic_vector(31 downto 0);
    signal iNsTr_62_2033 : std_logic_vector(31 downto 0);
    signal iNsTr_63_2039 : std_logic_vector(31 downto 0);
    signal iNsTr_64_2044 : std_logic_vector(31 downto 0);
    signal iNsTr_67_2818 : std_logic_vector(31 downto 0);
    signal iNsTr_68_2831 : std_logic_vector(31 downto 0);
    signal iNsTr_69_2836 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1727 : std_logic_vector(31 downto 0);
    signal iNsTr_70_2842 : std_logic_vector(31 downto 0);
    signal iNsTr_71_2848 : std_logic_vector(31 downto 0);
    signal iNsTr_72_2853 : std_logic_vector(31 downto 0);
    signal iNsTr_73_2859 : std_logic_vector(31 downto 0);
    signal iNsTr_74_2865 : std_logic_vector(0 downto 0);
    signal iNsTr_76_2419 : std_logic_vector(31 downto 0);
    signal iNsTr_77_2425 : std_logic_vector(31 downto 0);
    signal iNsTr_78_2431 : std_logic_vector(31 downto 0);
    signal iNsTr_79_2437 : std_logic_vector(31 downto 0);
    signal iNsTr_80_2443 : std_logic_vector(31 downto 0);
    signal iNsTr_81_2449 : std_logic_vector(31 downto 0);
    signal iNsTr_82_2455 : std_logic_vector(31 downto 0);
    signal iNsTr_83_2461 : std_logic_vector(31 downto 0);
    signal iNsTr_84_2467 : std_logic_vector(31 downto 0);
    signal iNsTr_85_2473 : std_logic_vector(31 downto 0);
    signal iNsTr_86_2478 : std_logic_vector(31 downto 0);
    signal iNsTr_87_2484 : std_logic_vector(31 downto 0);
    signal iNsTr_88_2489 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1730 : std_logic_vector(31 downto 0);
    signal iNsTr_92_2206 : std_logic_vector(31 downto 0);
    signal iNsTr_93_2212 : std_logic_vector(0 downto 0);
    signal iNsTr_94_2220 : std_logic_vector(0 downto 0);
    signal iNsTr_96_2904 : std_logic_vector(31 downto 0);
    signal iNsTr_97_2909 : std_logic_vector(31 downto 0);
    signal iNsTr_98_2915 : std_logic_vector(0 downto 0);
    signal indvarx_xnextx_xi_3220 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xix_xi19_2285 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xix_xi_2730 : std_logic_vector(31 downto 0);
    signal int_flux_err_temp_2x_x0_1669 : std_logic_vector(31 downto 0);
    signal int_flux_errx_x0_2888 : std_logic_vector(31 downto 0);
    signal int_speed_err_prevx_x0_1704 : std_logic_vector(31 downto 0);
    signal int_speed_errx_x0_1864 : std_logic_vector(31 downto 0);
    signal orx_xcond11x_xi_3160 : std_logic_vector(0 downto 0);
    signal orx_xcond11x_xix_xi15_2225 : std_logic_vector(0 downto 0);
    signal orx_xcond11x_xix_xi_2670 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xi_3214 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xix_xi18_2279 : std_logic_vector(0 downto 0);
    signal orx_xcondx_xix_xi_2724 : std_logic_vector(0 downto 0);
    signal phitmp31_3328 : std_logic_vector(31 downto 0);
    signal phitmp32_1917 : std_logic_vector(31 downto 0);
    signal phitmp33_3334 : std_logic_vector(31 downto 0);
    signal phitmp_3322 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xi_2990 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xix_xi4_2064 : std_logic_vector(31 downto 0);
    signal quotientx_x05x_xix_xix_xi_2509 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xi_3019 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xix_xi6_2092 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x03x_xix_xix_xi_2537 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xi_3069 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2141 : std_logic_vector(31 downto 0);
    signal shifted_divisorx_x0x_xlcssax_xix_xix_xi_2586 : std_logic_vector(31 downto 0);
    signal spd_lpf_prevx_x0_1697 : std_logic_vector(31 downto 0);
    signal speed_err_prevx_x0_1676 : std_logic_vector(31 downto 0);
    signal speed_refx_x0_1791 : std_logic_vector(31 downto 0);
    signal speed_refx_x1_1711 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xi_3177 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xix_xi17_2242 : std_logic_vector(31 downto 0);
    signal tempx_x012x_xix_xi_2687 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xi_3256 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xix_xi27_2332 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xlcssax_xix_xi_2777 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xphx_xix_xi14_2194 : std_logic_vector(31 downto 0);
    signal tempx_x0x_xphx_xix_xi_2639 : std_logic_vector(31 downto 0);
    signal theta_prevx_x0_1683 : std_logic_vector(31 downto 0);
    signal tmp10x_xi35_2963 : std_logic_vector(31 downto 0);
    signal tmp10x_xi35x_xin_2949 : std_logic_vector(31 downto 0);
    signal tmp10x_xix_xi1_1951 : std_logic_vector(31 downto 0);
    signal tmp10x_xix_xi_2400 : std_logic_vector(31 downto 0);
    signal tmp21x_xix_xi22_2313 : std_logic_vector(31 downto 0);
    signal tmp21x_xix_xi_2758 : std_logic_vector(31 downto 0);
    signal tmp25x_xi_3242 : std_logic_vector(31 downto 0);
    signal tmp25x_xix_xi23_2318 : std_logic_vector(31 downto 0);
    signal tmp25x_xix_xi_2763 : std_logic_vector(31 downto 0);
    signal tmp26x_xi_3247 : std_logic_vector(31 downto 0);
    signal tmp26x_xix_xi24_2323 : std_logic_vector(31 downto 0);
    signal tmp26x_xix_xi_2768 : std_logic_vector(31 downto 0);
    signal tmp3x_xi_3294 : std_logic_vector(31 downto 0);
    signal tmp3x_xix_xi28_2370 : std_logic_vector(31 downto 0);
    signal tmp3x_xix_xi_2815 : std_logic_vector(31 downto 0);
    signal tmp6x_xix_xi2_1955 : std_logic_vector(31 downto 0);
    signal torque_refx_x0_1920 : std_logic_vector(31 downto 0);
    signal type_cast_1666_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1668_wire : std_logic_vector(31 downto 0);
    signal type_cast_1673_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1675_wire : std_logic_vector(31 downto 0);
    signal type_cast_1680_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1682_wire : std_logic_vector(31 downto 0);
    signal type_cast_1687_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1689_wire : std_logic_vector(31 downto 0);
    signal type_cast_1694_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1696_wire : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1703_wire : std_logic_vector(31 downto 0);
    signal type_cast_1708_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1710_wire : std_logic_vector(31 downto 0);
    signal type_cast_1715_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1717_wire : std_logic_vector(31 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1782_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1794_wire : std_logic_vector(31 downto 0);
    signal type_cast_1796_wire : std_logic_vector(31 downto 0);
    signal type_cast_1798_wire : std_logic_vector(31 downto 0);
    signal type_cast_1803_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1824_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1839_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1867_wire : std_logic_vector(31 downto 0);
    signal type_cast_1870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1889_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1902_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1915_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1923_wire : std_logic_vector(31 downto 0);
    signal type_cast_1926_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1929_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1934_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1959_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1972_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1978_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1984_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1990_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1996_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2002_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2008_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2014_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2020_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2026_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2061_wire : std_logic_vector(31 downto 0);
    signal type_cast_2063_wire : std_logic_vector(31 downto 0);
    signal type_cast_2067_wire : std_logic_vector(31 downto 0);
    signal type_cast_2070_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2075_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2095_wire : std_logic_vector(31 downto 0);
    signal type_cast_2097_wire : std_logic_vector(31 downto 0);
    signal type_cast_2101_wire : std_logic_vector(31 downto 0);
    signal type_cast_2104_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2109_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2115_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2133_wire : std_logic_vector(31 downto 0);
    signal type_cast_2137_wire : std_logic_vector(31 downto 0);
    signal type_cast_2144_wire : std_logic_vector(31 downto 0);
    signal type_cast_2146_wire : std_logic_vector(31 downto 0);
    signal type_cast_2151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2153_wire : std_logic_vector(31 downto 0);
    signal type_cast_2180_wire : std_logic_vector(31 downto 0);
    signal type_cast_2188_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2190_wire : std_logic_vector(31 downto 0);
    signal type_cast_2197_wire : std_logic_vector(31 downto 0);
    signal type_cast_2199_wire : std_logic_vector(31 downto 0);
    signal type_cast_2204_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2215_wire : std_logic_vector(31 downto 0);
    signal type_cast_2218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2238_wire : std_logic_vector(31 downto 0);
    signal type_cast_2241_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2245_wire : std_logic_vector(31 downto 0);
    signal type_cast_2247_wire : std_logic_vector(31 downto 0);
    signal type_cast_2252_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2258_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2264_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2269_wire : std_logic_vector(31 downto 0);
    signal type_cast_2272_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2283_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2296_wire : std_logic_vector(31 downto 0);
    signal type_cast_2300_wire : std_logic_vector(31 downto 0);
    signal type_cast_2305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2311_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2329_wire : std_logic_vector(31 downto 0);
    signal type_cast_2331_wire : std_logic_vector(31 downto 0);
    signal type_cast_2335_wire : std_logic_vector(31 downto 0);
    signal type_cast_2337_wire : std_logic_vector(31 downto 0);
    signal type_cast_2342_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2348_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2354_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2376_wire : std_logic_vector(31 downto 0);
    signal type_cast_2379_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2389_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2404_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2435_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2453_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2459_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2465_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2471_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2506_wire : std_logic_vector(31 downto 0);
    signal type_cast_2508_wire : std_logic_vector(31 downto 0);
    signal type_cast_2512_wire : std_logic_vector(31 downto 0);
    signal type_cast_2515_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2520_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2540_wire : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire : std_logic_vector(31 downto 0);
    signal type_cast_2546_wire : std_logic_vector(31 downto 0);
    signal type_cast_2549_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2554_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2560_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2578_wire : std_logic_vector(31 downto 0);
    signal type_cast_2582_wire : std_logic_vector(31 downto 0);
    signal type_cast_2589_wire : std_logic_vector(31 downto 0);
    signal type_cast_2591_wire : std_logic_vector(31 downto 0);
    signal type_cast_2596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2598_wire : std_logic_vector(31 downto 0);
    signal type_cast_2625_wire : std_logic_vector(31 downto 0);
    signal type_cast_2633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2635_wire : std_logic_vector(31 downto 0);
    signal type_cast_2642_wire : std_logic_vector(31 downto 0);
    signal type_cast_2644_wire : std_logic_vector(31 downto 0);
    signal type_cast_2649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2655_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2660_wire : std_logic_vector(31 downto 0);
    signal type_cast_2663_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2683_wire : std_logic_vector(31 downto 0);
    signal type_cast_2686_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2690_wire : std_logic_vector(31 downto 0);
    signal type_cast_2692_wire : std_logic_vector(31 downto 0);
    signal type_cast_2697_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2709_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2714_wire : std_logic_vector(31 downto 0);
    signal type_cast_2717_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2728_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2741_wire : std_logic_vector(31 downto 0);
    signal type_cast_2745_wire : std_logic_vector(31 downto 0);
    signal type_cast_2750_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2756_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2774_wire : std_logic_vector(31 downto 0);
    signal type_cast_2776_wire : std_logic_vector(31 downto 0);
    signal type_cast_2780_wire : std_logic_vector(31 downto 0);
    signal type_cast_2782_wire : std_logic_vector(31 downto 0);
    signal type_cast_2787_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2793_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2799_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2821_wire : std_logic_vector(31 downto 0);
    signal type_cast_2824_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2829_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2839_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2846_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2857_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2876_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2891_wire : std_logic_vector(31 downto 0);
    signal type_cast_2894_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2897_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2902_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2913_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2926_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2939_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2952_wire : std_logic_vector(31 downto 0);
    signal type_cast_2955_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2958_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2967_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2973_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2979_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2987_wire : std_logic_vector(31 downto 0);
    signal type_cast_2989_wire : std_logic_vector(31 downto 0);
    signal type_cast_2993_wire : std_logic_vector(31 downto 0);
    signal type_cast_2996_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3001_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3007_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3022_wire : std_logic_vector(31 downto 0);
    signal type_cast_3025_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3029_wire : std_logic_vector(31 downto 0);
    signal type_cast_3032_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3043_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3061_wire : std_logic_vector(31 downto 0);
    signal type_cast_3065_wire : std_logic_vector(31 downto 0);
    signal type_cast_3073_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3075_wire : std_logic_vector(31 downto 0);
    signal type_cast_3080_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3082_wire : std_logic_vector(31 downto 0);
    signal type_cast_3097_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3110_wire : std_logic_vector(31 downto 0);
    signal type_cast_3115_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3121_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3127_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3139_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3145_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3150_wire : std_logic_vector(31 downto 0);
    signal type_cast_3153_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3173_wire : std_logic_vector(31 downto 0);
    signal type_cast_3176_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3180_wire : std_logic_vector(31 downto 0);
    signal type_cast_3182_wire : std_logic_vector(31 downto 0);
    signal type_cast_3187_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3199_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3204_wire : std_logic_vector(31 downto 0);
    signal type_cast_3207_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3231_wire : std_logic_vector(31 downto 0);
    signal type_cast_3235_wire : std_logic_vector(31 downto 0);
    signal type_cast_3240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3253_wire : std_logic_vector(31 downto 0);
    signal type_cast_3255_wire : std_logic_vector(31 downto 0);
    signal type_cast_3259_wire : std_logic_vector(31 downto 0);
    signal type_cast_3261_wire : std_logic_vector(31 downto 0);
    signal type_cast_3266_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3272_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3278_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3300_wire : std_logic_vector(31 downto 0);
    signal type_cast_3303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3320_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3326_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3332_wire_constant : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xi_2984 : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xix_xi3_2058 : std_logic_vector(31 downto 0);
    signal xx_x016x_xix_xix_xi_2503 : std_logic_vector(31 downto 0);
    signal xx_x0x_xix_xix_xi12_2184 : std_logic_vector(31 downto 0);
    signal xx_x0x_xix_xix_xi_2629 : std_logic_vector(31 downto 0);
    signal xx_xlcssa10_2297 : std_logic_vector(31 downto 0);
    signal xx_xlcssa11_2293 : std_logic_vector(31 downto 0);
    signal xx_xlcssa12_2134 : std_logic_vector(31 downto 0);
    signal xx_xlcssa13_2130 : std_logic_vector(31 downto 0);
    signal xx_xlcssa14_2177 : std_logic_vector(31 downto 0);
    signal xx_xlcssa1_3228 : std_logic_vector(31 downto 0);
    signal xx_xlcssa2_3062 : std_logic_vector(31 downto 0);
    signal xx_xlcssa3_3058 : std_logic_vector(31 downto 0);
    signal xx_xlcssa4_3107 : std_logic_vector(31 downto 0);
    signal xx_xlcssa5_2742 : std_logic_vector(31 downto 0);
    signal xx_xlcssa6_2738 : std_logic_vector(31 downto 0);
    signal xx_xlcssa7_2579 : std_logic_vector(31 downto 0);
    signal xx_xlcssa8_2575 : std_logic_vector(31 downto 0);
    signal xx_xlcssa9_2622 : std_logic_vector(31 downto 0);
    signal xx_xlcssa_3232 : std_logic_vector(31 downto 0);
    signal xx_xnotx_xi21_2307 : std_logic_vector(31 downto 0);
    signal xx_xnotx_xi_2752 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    expr_2047_wire_constant <= "00000000000000000000000000000000";
    expr_2050_wire_constant <= "00000000000000000000000000000001";
    expr_2492_wire_constant <= "00000000000000000000000000000000";
    expr_2495_wire_constant <= "00000000000000000000000000000001";
    type_cast_1666_wire_constant <= "00000000000000000000000000000000";
    type_cast_1673_wire_constant <= "00000000000000000000000000000000";
    type_cast_1680_wire_constant <= "00000000000000000000000000000000";
    type_cast_1687_wire_constant <= "00000000000000000000000000000000";
    type_cast_1694_wire_constant <= "00000000000000000000000000000000";
    type_cast_1701_wire_constant <= "00000000000000000000000000000000";
    type_cast_1708_wire_constant <= "00000000000000000000000000000000";
    type_cast_1715_wire_constant <= "00000000000000000000000000000000";
    type_cast_1754_wire_constant <= "0011111110101001100110011001100110011001100110011001100110011010";
    type_cast_1782_wire_constant <= "1011111110101001100110011001100110011001100110011001100110011010";
    type_cast_1803_wire_constant <= "00111111001100110011001100110011";
    type_cast_1824_wire_constant <= "00111001100000110001001001101111";
    type_cast_1839_wire_constant <= "1100000000100100000000000000000000000000000000000000000000000000";
    type_cast_1852_wire_constant <= "0100000000100100000000000000000000000000000000000000000000000000";
    type_cast_1870_wire_constant <= "11000001001000000000000000000000";
    type_cast_1873_wire_constant <= "01000001001000000000000000000000";
    type_cast_1878_wire_constant <= "01000000101000000000000000000000";
    type_cast_1889_wire_constant <= "11000001101000000000000000000000";
    type_cast_1902_wire_constant <= "01000001101000000000000000000000";
    type_cast_1915_wire_constant <= "00111110101100010111000110101010";
    type_cast_1926_wire_constant <= "11000000110111011100111000010100";
    type_cast_1929_wire_constant <= "01000000110111011100111000010100";
    type_cast_1934_wire_constant <= "00111001110010111011111000010101";
    type_cast_1945_wire_constant <= "01000000111110010100110011010001";
    type_cast_1959_wire_constant <= "00000000000000000000000000000000";
    type_cast_1972_wire_constant <= "00000000000000000000000000010111";
    type_cast_1978_wire_constant <= "00000000000000000000000011111111";
    type_cast_1984_wire_constant <= "00000000000000000000000000010111";
    type_cast_1990_wire_constant <= "00000000000000000000000011111111";
    type_cast_1996_wire_constant <= "00000000000000000000000000000111";
    type_cast_2002_wire_constant <= "00111111111111111111111110000000";
    type_cast_2008_wire_constant <= "01000000000000000000000000000000";
    type_cast_2014_wire_constant <= "00000000000000000000000000000111";
    type_cast_2020_wire_constant <= "00000000000000001111111111111111";
    type_cast_2026_wire_constant <= "00000000000000010000000000000000";
    type_cast_2037_wire_constant <= "10000000000000000000000000000000";
    type_cast_2070_wire_constant <= "00000000000000000000000000000000";
    type_cast_2075_wire_constant <= "00000000000000000000000000000001";
    type_cast_2104_wire_constant <= "00000000000000000000000000000001";
    type_cast_2109_wire_constant <= "00000000000000000000000000000001";
    type_cast_2115_wire_constant <= "00000000000000000000000000000001";
    type_cast_2151_wire_constant <= "00000000000000000000000000000001";
    type_cast_2188_wire_constant <= "11111111111111111111111111111111";
    type_cast_2204_wire_constant <= "00000000100000000000000000000000";
    type_cast_2210_wire_constant <= "00000000000000000000000000000000";
    type_cast_2218_wire_constant <= "00000000000000000000000000000000";
    type_cast_2241_wire_constant <= "00000000000000000000000000000000";
    type_cast_2252_wire_constant <= "00000000000000000000000000000001";
    type_cast_2258_wire_constant <= "00000000100000000000000000000000";
    type_cast_2264_wire_constant <= "00000000000000000000000000000000";
    type_cast_2272_wire_constant <= "00000000000000000000000000000000";
    type_cast_2283_wire_constant <= "00000000000000000000000000000001";
    type_cast_2305_wire_constant <= "11111111111111111111111100000000";
    type_cast_2311_wire_constant <= "00000000000000000000000011111111";
    type_cast_2342_wire_constant <= "00000000011111111111111111111111";
    type_cast_2348_wire_constant <= "00000000000000000000000000010111";
    type_cast_2354_wire_constant <= "01000100000000000000000000000000";
    type_cast_2379_wire_constant <= "00000000000000000000000000000000";
    type_cast_2389_wire_constant <= "00111000010100011011011100010111";
    type_cast_2404_wire_constant <= "00000000000000000000000000000000";
    type_cast_2417_wire_constant <= "00000000000000000000000000010111";
    type_cast_2423_wire_constant <= "00000000000000000000000011111111";
    type_cast_2429_wire_constant <= "00000000000000000000000000010111";
    type_cast_2435_wire_constant <= "00000000000000000000000011111111";
    type_cast_2441_wire_constant <= "00000000000000000000000000000111";
    type_cast_2447_wire_constant <= "00111111111111111111111110000000";
    type_cast_2453_wire_constant <= "01000000000000000000000000000000";
    type_cast_2459_wire_constant <= "00000000000000000000000000000111";
    type_cast_2465_wire_constant <= "00000000000000001111111111111111";
    type_cast_2471_wire_constant <= "00000000000000010000000000000000";
    type_cast_2482_wire_constant <= "10000000000000000000000000000000";
    type_cast_2515_wire_constant <= "00000000000000000000000000000000";
    type_cast_2520_wire_constant <= "00000000000000000000000000000001";
    type_cast_2549_wire_constant <= "00000000000000000000000000000001";
    type_cast_2554_wire_constant <= "00000000000000000000000000000001";
    type_cast_2560_wire_constant <= "00000000000000000000000000000001";
    type_cast_2596_wire_constant <= "00000000000000000000000000000001";
    type_cast_2633_wire_constant <= "11111111111111111111111111111111";
    type_cast_2649_wire_constant <= "00000000100000000000000000000000";
    type_cast_2655_wire_constant <= "00000000000000000000000000000000";
    type_cast_2663_wire_constant <= "00000000000000000000000000000000";
    type_cast_2686_wire_constant <= "00000000000000000000000000000000";
    type_cast_2697_wire_constant <= "00000000000000000000000000000001";
    type_cast_2703_wire_constant <= "00000000100000000000000000000000";
    type_cast_2709_wire_constant <= "00000000000000000000000000000000";
    type_cast_2717_wire_constant <= "00000000000000000000000000000000";
    type_cast_2728_wire_constant <= "00000000000000000000000000000001";
    type_cast_2750_wire_constant <= "11111111111111111111111100000000";
    type_cast_2756_wire_constant <= "00000000000000000000000011111111";
    type_cast_2787_wire_constant <= "00000000011111111111111111111111";
    type_cast_2793_wire_constant <= "00000000000000000000000000010111";
    type_cast_2799_wire_constant <= "01000100000000000000000000000000";
    type_cast_2824_wire_constant <= "00000000000000000000000000000000";
    type_cast_2829_wire_constant <= "00111011101001000100110001111011";
    type_cast_2839_wire_constant <= "00111110100110011001100110011010";
    type_cast_2846_wire_constant <= "00111000010100011011011100010111";
    type_cast_2857_wire_constant <= "01000010010010000000000000000000";
    type_cast_2863_wire_constant <= "10111111100000000000000000000000";
    type_cast_2876_wire_constant <= "00111111100000000000000000000000";
    type_cast_2894_wire_constant <= "10111111100000000000000000000000";
    type_cast_2897_wire_constant <= "00111111100000000000000000000000";
    type_cast_2902_wire_constant <= "01000010001000000000000000000000";
    type_cast_2913_wire_constant <= "11000000000000000000000000000000";
    type_cast_2926_wire_constant <= "01000000000000000000000000000000";
    type_cast_2939_wire_constant <= "00000000000000000000000000000000";
    type_cast_2955_wire_constant <= "11000000000000000000000000000000";
    type_cast_2958_wire_constant <= "01000000000000000000000000000000";
    type_cast_2967_wire_constant <= "00000000000000000000000000000111";
    type_cast_2973_wire_constant <= "00111111111111111111111110000000";
    type_cast_2979_wire_constant <= "01000000000000000000000000000000";
    type_cast_2996_wire_constant <= "00000000000000000000000000000000";
    type_cast_3001_wire_constant <= "00000000000000000000000000000001";
    type_cast_3007_wire_constant <= "00000000000000011001111010000011";
    type_cast_3025_wire_constant <= "00000000000000011001111010000011";
    type_cast_3032_wire_constant <= "00000000000000000000000000000001";
    type_cast_3037_wire_constant <= "00000000000000000000000000000001";
    type_cast_3043_wire_constant <= "00000000000000000000000000000001";
    type_cast_3073_wire_constant <= "00000000000000011001111010000011";
    type_cast_3080_wire_constant <= "00000000000000000000000000000001";
    type_cast_3097_wire_constant <= "00000000000000011001111010000011";
    type_cast_3115_wire_constant <= "00000000000000000000000000010111";
    type_cast_3121_wire_constant <= "10000000000000000000000000000000";
    type_cast_3127_wire_constant <= "00000000000000000000000011111111";
    type_cast_3133_wire_constant <= "11111111111111111111111110000010";
    type_cast_3139_wire_constant <= "00000000100000000000000000000000";
    type_cast_3145_wire_constant <= "00000000000000000000000000000000";
    type_cast_3153_wire_constant <= "00000000000000000000000000000000";
    type_cast_3176_wire_constant <= "00000000000000000000000000000000";
    type_cast_3187_wire_constant <= "00000000000000000000000000000001";
    type_cast_3193_wire_constant <= "00000000100000000000000000000000";
    type_cast_3199_wire_constant <= "00000000000000000000000000000000";
    type_cast_3207_wire_constant <= "00000000000000000000000000000000";
    type_cast_3218_wire_constant <= "00000000000000000000000000000001";
    type_cast_3240_wire_constant <= "11111111111111111111111110000001";
    type_cast_3266_wire_constant <= "00000000011111111111111111111111";
    type_cast_3272_wire_constant <= "00000000000000000000000000010111";
    type_cast_3278_wire_constant <= "01000100000000000000000000000000";
    type_cast_3303_wire_constant <= "00000000000000000000000000000000";
    type_cast_3320_wire_constant <= "00111110100110011001100110011010";
    type_cast_3326_wire_constant <= "00111111011111111110000010001011";
    type_cast_3332_wire_constant <= "00111111011111101011011101100111";
    phi_stmt_1662: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1666_wire_constant & type_cast_1668_wire;
      req <= phi_stmt_1662_req_0 & phi_stmt_1662_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1662_ack_0,
          idata => idata,
          odata => flux_rotor_lpf_prevx_x0_1662,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1662
    phi_stmt_1669: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1673_wire_constant & type_cast_1675_wire;
      req <= phi_stmt_1669_req_0 & phi_stmt_1669_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1669_ack_0,
          idata => idata,
          odata => int_flux_err_temp_2x_x0_1669,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1669
    phi_stmt_1676: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1680_wire_constant & type_cast_1682_wire;
      req <= phi_stmt_1676_req_0 & phi_stmt_1676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1676_ack_0,
          idata => idata,
          odata => speed_err_prevx_x0_1676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1676
    phi_stmt_1683: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1687_wire_constant & type_cast_1689_wire;
      req <= phi_stmt_1683_req_0 & phi_stmt_1683_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1683_ack_0,
          idata => idata,
          odata => theta_prevx_x0_1683,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1683
    phi_stmt_1690: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1694_wire_constant & type_cast_1696_wire;
      req <= phi_stmt_1690_req_0 & phi_stmt_1690_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1690_ack_0,
          idata => idata,
          odata => flux_rotor_prevx_x0_1690,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1690
    phi_stmt_1697: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1701_wire_constant & type_cast_1703_wire;
      req <= phi_stmt_1697_req_0 & phi_stmt_1697_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1697_ack_0,
          idata => idata,
          odata => spd_lpf_prevx_x0_1697,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1697
    phi_stmt_1704: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1708_wire_constant & type_cast_1710_wire;
      req <= phi_stmt_1704_req_0 & phi_stmt_1704_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1704_ack_0,
          idata => idata,
          odata => int_speed_err_prevx_x0_1704,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1704
    phi_stmt_1711: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1715_wire_constant & type_cast_1717_wire;
      req <= phi_stmt_1711_req_0 & phi_stmt_1711_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1711_ack_0,
          idata => idata,
          odata => speed_refx_x1_1711,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1711
    phi_stmt_1791: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1794_wire & type_cast_1796_wire & type_cast_1798_wire;
      req <= phi_stmt_1791_req_0 & phi_stmt_1791_req_1 & phi_stmt_1791_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1791_ack_0,
          idata => idata,
          odata => speed_refx_x0_1791,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1791
    phi_stmt_1864: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1867_wire & type_cast_1870_wire_constant & type_cast_1873_wire_constant;
      req <= phi_stmt_1864_req_0 & phi_stmt_1864_req_1 & phi_stmt_1864_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1864_ack_0,
          idata => idata,
          odata => int_speed_errx_x0_1864,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1864
    phi_stmt_1920: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1923_wire & type_cast_1926_wire_constant & type_cast_1929_wire_constant;
      req <= phi_stmt_1920_req_0 & phi_stmt_1920_req_1 & phi_stmt_1920_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1920_ack_0,
          idata => idata,
          odata => torque_refx_x0_1920,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1920
    phi_stmt_2058: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2061_wire & type_cast_2063_wire;
      req <= phi_stmt_2058_req_0 & phi_stmt_2058_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2058_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xix_xi3_2058,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2058
    phi_stmt_2064: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2067_wire & type_cast_2070_wire_constant;
      req <= phi_stmt_2064_req_0 & phi_stmt_2064_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2064_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xix_xi4_2064,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2064
    phi_stmt_2092: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2095_wire & type_cast_2097_wire;
      req <= phi_stmt_2092_req_0 & phi_stmt_2092_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2092_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xix_xi6_2092,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2092
    phi_stmt_2098: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2101_wire & type_cast_2104_wire_constant;
      req <= phi_stmt_2098_req_0 & phi_stmt_2098_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2098_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xix_xi7_2098,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2098
    phi_stmt_2130: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2133_wire;
      req(0) <= phi_stmt_2130_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2130_ack_0,
          idata => idata,
          odata => xx_xlcssa13_2130,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2130
    phi_stmt_2134: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2137_wire;
      req(0) <= phi_stmt_2134_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2134_ack_0,
          idata => idata,
          odata => xx_xlcssa12_2134,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2134
    phi_stmt_2141: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2144_wire & type_cast_2146_wire;
      req <= phi_stmt_2141_req_0 & phi_stmt_2141_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2141_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2141,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2141
    phi_stmt_2147: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2151_wire_constant & type_cast_2153_wire;
      req <= phi_stmt_2147_req_0 & phi_stmt_2147_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2147_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xix_xi10_2147,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2147
    phi_stmt_2177: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2180_wire;
      req(0) <= phi_stmt_2177_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2177_ack_0,
          idata => idata,
          odata => xx_xlcssa14_2177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2177
    phi_stmt_2184: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2188_wire_constant & type_cast_2190_wire;
      req <= phi_stmt_2184_req_0 & phi_stmt_2184_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2184_ack_0,
          idata => idata,
          odata => xx_x0x_xix_xix_xi12_2184,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2184
    phi_stmt_2194: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2197_wire & type_cast_2199_wire;
      req <= phi_stmt_2194_req_0 & phi_stmt_2194_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2194_ack_0,
          idata => idata,
          odata => tempx_x0x_xphx_xix_xi14_2194,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2194
    phi_stmt_2235: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2238_wire & type_cast_2241_wire_constant;
      req <= phi_stmt_2235_req_0 & phi_stmt_2235_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2235_ack_0,
          idata => idata,
          odata => iNsTr_140_2235,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2235
    phi_stmt_2242: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2245_wire & type_cast_2247_wire;
      req <= phi_stmt_2242_req_0 & phi_stmt_2242_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2242_ack_0,
          idata => idata,
          odata => tempx_x012x_xix_xi17_2242,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2242
    phi_stmt_2293: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2296_wire;
      req(0) <= phi_stmt_2293_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2293_ack_0,
          idata => idata,
          odata => xx_xlcssa11_2293,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2293
    phi_stmt_2297: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2300_wire;
      req(0) <= phi_stmt_2297_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2297_ack_0,
          idata => idata,
          odata => xx_xlcssa10_2297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2297
    phi_stmt_2326: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2329_wire & type_cast_2331_wire;
      req <= phi_stmt_2326_req_0 & phi_stmt_2326_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2326_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xix_xi26_2326,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2326
    phi_stmt_2332: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2335_wire & type_cast_2337_wire;
      req <= phi_stmt_2332_req_0 & phi_stmt_2332_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2332_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xix_xi27_2332,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2332
    phi_stmt_2373: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2376_wire & type_cast_2379_wire_constant;
      req <= phi_stmt_2373_req_0 & phi_stmt_2373_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2373_ack_0,
          idata => idata,
          odata => iNsTr_46_2373,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2373
    phi_stmt_2503: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2506_wire & type_cast_2508_wire;
      req <= phi_stmt_2503_req_0 & phi_stmt_2503_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2503_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xix_xi_2503,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2503
    phi_stmt_2509: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2512_wire & type_cast_2515_wire_constant;
      req <= phi_stmt_2509_req_0 & phi_stmt_2509_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2509_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xix_xi_2509,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2509
    phi_stmt_2537: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2540_wire & type_cast_2542_wire;
      req <= phi_stmt_2537_req_0 & phi_stmt_2537_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2537_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xix_xi_2537,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2537
    phi_stmt_2543: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2546_wire & type_cast_2549_wire_constant;
      req <= phi_stmt_2543_req_0 & phi_stmt_2543_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2543_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xix_xi_2543,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2543
    phi_stmt_2575: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2578_wire;
      req(0) <= phi_stmt_2575_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2575_ack_0,
          idata => idata,
          odata => xx_xlcssa8_2575,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2575
    phi_stmt_2579: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2582_wire;
      req(0) <= phi_stmt_2579_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2579_ack_0,
          idata => idata,
          odata => xx_xlcssa7_2579,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2579
    phi_stmt_2586: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2589_wire & type_cast_2591_wire;
      req <= phi_stmt_2586_req_0 & phi_stmt_2586_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2586_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xix_xi_2586,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2586
    phi_stmt_2592: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2596_wire_constant & type_cast_2598_wire;
      req <= phi_stmt_2592_req_0 & phi_stmt_2592_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2592_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xix_xi_2592,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2592
    phi_stmt_2622: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2625_wire;
      req(0) <= phi_stmt_2622_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2622_ack_0,
          idata => idata,
          odata => xx_xlcssa9_2622,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2622
    phi_stmt_2629: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2633_wire_constant & type_cast_2635_wire;
      req <= phi_stmt_2629_req_0 & phi_stmt_2629_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2629_ack_0,
          idata => idata,
          odata => xx_x0x_xix_xix_xi_2629,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2629
    phi_stmt_2639: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2642_wire & type_cast_2644_wire;
      req <= phi_stmt_2639_req_0 & phi_stmt_2639_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2639_ack_0,
          idata => idata,
          odata => tempx_x0x_xphx_xix_xi_2639,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2639
    phi_stmt_2680: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2683_wire & type_cast_2686_wire_constant;
      req <= phi_stmt_2680_req_0 & phi_stmt_2680_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2680_ack_0,
          idata => idata,
          odata => iNsTr_156_2680,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2680
    phi_stmt_2687: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2690_wire & type_cast_2692_wire;
      req <= phi_stmt_2687_req_0 & phi_stmt_2687_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2687_ack_0,
          idata => idata,
          odata => tempx_x012x_xix_xi_2687,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2687
    phi_stmt_2738: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2741_wire;
      req(0) <= phi_stmt_2738_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2738_ack_0,
          idata => idata,
          odata => xx_xlcssa6_2738,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2738
    phi_stmt_2742: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2745_wire;
      req(0) <= phi_stmt_2742_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2742_ack_0,
          idata => idata,
          odata => xx_xlcssa5_2742,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2742
    phi_stmt_2771: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2774_wire & type_cast_2776_wire;
      req <= phi_stmt_2771_req_0 & phi_stmt_2771_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2771_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xix_xi_2771,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2771
    phi_stmt_2777: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2780_wire & type_cast_2782_wire;
      req <= phi_stmt_2777_req_0 & phi_stmt_2777_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2777_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xix_xi_2777,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2777
    phi_stmt_2818: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2821_wire & type_cast_2824_wire_constant;
      req <= phi_stmt_2818_req_0 & phi_stmt_2818_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2818_ack_0,
          idata => idata,
          odata => iNsTr_67_2818,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2818
    phi_stmt_2888: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2891_wire & type_cast_2894_wire_constant & type_cast_2897_wire_constant;
      req <= phi_stmt_2888_req_0 & phi_stmt_2888_req_1 & phi_stmt_2888_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2888_ack_0,
          idata => idata,
          odata => int_flux_errx_x0_2888,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2888
    phi_stmt_2949: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2952_wire & type_cast_2955_wire_constant & type_cast_2958_wire_constant;
      req <= phi_stmt_2949_req_0 & phi_stmt_2949_req_1 & phi_stmt_2949_req_2;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 3,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2949_ack_0,
          idata => idata,
          odata => tmp10x_xi35x_xin_2949,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2949
    phi_stmt_2984: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2987_wire & type_cast_2989_wire;
      req <= phi_stmt_2984_req_0 & phi_stmt_2984_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2984_ack_0,
          idata => idata,
          odata => xx_x016x_xix_xi_2984,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2984
    phi_stmt_2990: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2993_wire & type_cast_2996_wire_constant;
      req <= phi_stmt_2990_req_0 & phi_stmt_2990_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2990_ack_0,
          idata => idata,
          odata => quotientx_x05x_xix_xi_2990,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2990
    phi_stmt_3019: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3022_wire & type_cast_3025_wire_constant;
      req <= phi_stmt_3019_req_0 & phi_stmt_3019_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3019_ack_0,
          idata => idata,
          odata => shifted_divisorx_x03x_xix_xi_3019,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3019
    phi_stmt_3026: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3029_wire & type_cast_3032_wire_constant;
      req <= phi_stmt_3026_req_0 & phi_stmt_3026_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3026_ack_0,
          idata => idata,
          odata => curr_quotientx_x02x_xix_xi_3026,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3026
    phi_stmt_3058: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3061_wire;
      req(0) <= phi_stmt_3058_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3058_ack_0,
          idata => idata,
          odata => xx_xlcssa3_3058,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3058
    phi_stmt_3062: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3065_wire;
      req(0) <= phi_stmt_3062_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3062_ack_0,
          idata => idata,
          odata => xx_xlcssa2_3062,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3062
    phi_stmt_3069: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3073_wire_constant & type_cast_3075_wire;
      req <= phi_stmt_3069_req_0 & phi_stmt_3069_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3069_ack_0,
          idata => idata,
          odata => shifted_divisorx_x0x_xlcssax_xix_xi_3069,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3069
    phi_stmt_3076: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3080_wire_constant & type_cast_3082_wire;
      req <= phi_stmt_3076_req_0 & phi_stmt_3076_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3076_ack_0,
          idata => idata,
          odata => curr_quotientx_x0x_xlcssax_xix_xi_3076,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3076
    phi_stmt_3107: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3110_wire;
      req(0) <= phi_stmt_3107_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3107_ack_0,
          idata => idata,
          odata => xx_xlcssa4_3107,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3107
    phi_stmt_3170: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3173_wire & type_cast_3176_wire_constant;
      req <= phi_stmt_3170_req_0 & phi_stmt_3170_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3170_ack_0,
          idata => idata,
          odata => iNsTr_211_3170,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3170
    phi_stmt_3177: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3180_wire & type_cast_3182_wire;
      req <= phi_stmt_3177_req_0 & phi_stmt_3177_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3177_ack_0,
          idata => idata,
          odata => tempx_x012x_xi_3177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3177
    phi_stmt_3228: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3231_wire;
      req(0) <= phi_stmt_3228_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3228_ack_0,
          idata => idata,
          odata => xx_xlcssa1_3228,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3228
    phi_stmt_3232: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3235_wire;
      req(0) <= phi_stmt_3232_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3232_ack_0,
          idata => idata,
          odata => xx_xlcssa_3232,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3232
    phi_stmt_3250: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3253_wire & type_cast_3255_wire;
      req <= phi_stmt_3250_req_0 & phi_stmt_3250_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3250_ack_0,
          idata => idata,
          odata => expx_x0x_xlcssax_xi_3250,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3250
    phi_stmt_3256: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3259_wire & type_cast_3261_wire;
      req <= phi_stmt_3256_req_0 & phi_stmt_3256_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3256_ack_0,
          idata => idata,
          odata => tempx_x0x_xlcssax_xi_3256,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3256
    phi_stmt_3297: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3300_wire & type_cast_3303_wire_constant;
      req <= phi_stmt_3297_req_0 & phi_stmt_3297_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3297_ack_0,
          idata => idata,
          odata => iNsTr_173_3297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3297
    type_cast_1668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1668_inst_req_0;
      type_cast_1668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1668_inst_req_1;
      type_cast_1668_inst_ack_1<= rack(0);
      type_cast_1668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1668_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp33_3334,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1668_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1675_inst_req_0;
      type_cast_1675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1675_inst_req_1;
      type_cast_1675_inst_ack_1<= rack(0);
      type_cast_1675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1675_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_72_2853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1675_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1682_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1682_inst_req_0;
      type_cast_1682_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1682_inst_req_1;
      type_cast_1682_inst_ack_1<= rack(0);
      type_cast_1682_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1682_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_21_1815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1682_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1689_inst_req_0;
      type_cast_1689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1689_inst_req_1;
      type_cast_1689_inst_ack_1<= rack(0);
      type_cast_1689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1689_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_49_2396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1689_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1696_inst_req_0;
      type_cast_1696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1696_inst_req_1;
      type_cast_1696_inst_ack_1<= rack(0);
      type_cast_1696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1696_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp31_3328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1696_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1703_inst_req_0;
      type_cast_1703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1703_inst_req_1;
      type_cast_1703_inst_ack_1<= rack(0);
      type_cast_1703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1703_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_3322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1703_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1710_inst_req_0;
      type_cast_1710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1710_inst_req_1;
      type_cast_1710_inst_ack_1<= rack(0);
      type_cast_1710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1710_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_24_1831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1710_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1717_inst_req_0;
      type_cast_1717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1717_inst_req_1;
      type_cast_1717_inst_ack_1<= rack(0);
      type_cast_1717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1717_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => speed_refx_x0_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1717_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1794_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1794_inst_req_0;
      type_cast_1794_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1794_inst_req_1;
      type_cast_1794_inst_ack_1<= rack(0);
      type_cast_1794_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1794_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_15_1760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1794_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1796_inst_req_0;
      type_cast_1796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1796_inst_req_1;
      type_cast_1796_inst_ack_1<= rack(0);
      type_cast_1796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1796_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_30_1788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1796_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1798_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1798_inst_req_0;
      type_cast_1798_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1798_inst_req_1;
      type_cast_1798_inst_ack_1<= rack(0);
      type_cast_1798_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1798_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => speed_refx_x1_1711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1798_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1867_inst_req_0;
      type_cast_1867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1867_inst_req_1;
      type_cast_1867_inst_ack_1<= rack(0);
      type_cast_1867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1867_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_24_1831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1867_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1923_inst_req_0;
      type_cast_1923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1923_inst_req_1;
      type_cast_1923_inst_ack_1<= rack(0);
      type_cast_1923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1923_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp32_1917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1950_inst_req_0;
      type_cast_1950_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1950_inst_req_1;
      type_cast_1950_inst_ack_1<= rack(0);
      type_cast_1950_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1950_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_40_1947,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xix_xi1_1951,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1954_inst_req_0;
      type_cast_1954_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1954_inst_req_1;
      type_cast_1954_inst_ack_1<= rack(0);
      type_cast_1954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1954_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_39_1941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6x_xix_xi2_1955,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_137_2164,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2063_inst_req_0;
      type_cast_2063_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2063_inst_req_1;
      type_cast_2063_inst_ack_1<= rack(0);
      type_cast_2063_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2063_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_58_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2063_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2067_inst_req_0;
      type_cast_2067_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2067_inst_req_1;
      type_cast_2067_inst_ack_1<= rack(0);
      type_cast_2067_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2067_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_136_2159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2067_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2095_inst_req_0;
      type_cast_2095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2095_inst_req_1;
      type_cast_2095_inst_ack_1<= rack(0);
      type_cast_2095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2095_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_162_2111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2095_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2097_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2097_inst_req_0;
      type_cast_2097_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2097_inst_req_1;
      type_cast_2097_inst_ack_1<= rack(0);
      type_cast_2097_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2097_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_61_2028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2097_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2101_inst_req_0;
      type_cast_2101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2101_inst_req_1;
      type_cast_2101_inst_ack_1<= rack(0);
      type_cast_2101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2101_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_163_2117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2101_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2133_inst_req_0;
      type_cast_2133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2133_inst_req_1;
      type_cast_2133_inst_ack_1<= rack(0);
      type_cast_2133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2133_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_163_2117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2133_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2137_inst_req_0;
      type_cast_2137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2137_inst_req_1;
      type_cast_2137_inst_ack_1<= rack(0);
      type_cast_2137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2137_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_162_2111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2137_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2144_inst_req_0;
      type_cast_2144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2144_inst_req_1;
      type_cast_2144_inst_ack_1<= rack(0);
      type_cast_2144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2144_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_61_2028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2144_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2146_inst_req_0;
      type_cast_2146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2146_inst_req_1;
      type_cast_2146_inst_ack_1<= rack(0);
      type_cast_2146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2146_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa12_2134,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2146_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2153_inst_req_0;
      type_cast_2153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2153_inst_req_1;
      type_cast_2153_inst_ack_1<= rack(0);
      type_cast_2153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2153_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa13_2130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_136_2159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2180_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2190_inst_req_0;
      type_cast_2190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2190_inst_req_1;
      type_cast_2190_inst_ack_1<= rack(0);
      type_cast_2190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2190_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa14_2177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2190_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2197_inst_req_0;
      type_cast_2197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2197_inst_req_1;
      type_cast_2197_inst_ack_1<= rack(0);
      type_cast_2197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2197_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_x0x_xix_xix_xi12_2184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2197_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_58_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2238_inst_req_0;
      type_cast_2238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2238_inst_req_1;
      type_cast_2238_inst_ack_1<= rack(0);
      type_cast_2238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2238_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xix_xi19_2285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2238_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2245_inst_req_0;
      type_cast_2245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2245_inst_req_1;
      type_cast_2245_inst_ack_1<= rack(0);
      type_cast_2245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2245_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_141_2254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2245_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2247_inst_req_0;
      type_cast_2247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2247_inst_req_1;
      type_cast_2247_inst_ack_1<= rack(0);
      type_cast_2247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2247_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi14_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2247_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2296_inst_req_0;
      type_cast_2296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2296_inst_req_1;
      type_cast_2296_inst_ack_1<= rack(0);
      type_cast_2296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2296_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_141_2254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2296_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2300_inst_req_0;
      type_cast_2300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2300_inst_req_1;
      type_cast_2300_inst_ack_1<= rack(0);
      type_cast_2300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2300_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_140_2235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2300_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2329_inst_req_0;
      type_cast_2329_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2329_inst_req_1;
      type_cast_2329_inst_ack_1<= rack(0);
      type_cast_2329_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2329_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xix_xi24_2323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2329_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2331_inst_req_0;
      type_cast_2331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2331_inst_req_1;
      type_cast_2331_inst_ack_1<= rack(0);
      type_cast_2331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2331_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_64_2044,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2331_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2335_inst_req_0;
      type_cast_2335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2335_inst_req_1;
      type_cast_2335_inst_ack_1<= rack(0);
      type_cast_2335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2335_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa11_2293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2335_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2337_inst_req_0;
      type_cast_2337_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2337_inst_req_1;
      type_cast_2337_inst_ack_1<= rack(0);
      type_cast_2337_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2337_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi14_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2337_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2369_inst_req_0;
      type_cast_2369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2369_inst_req_1;
      type_cast_2369_inst_ack_1<= rack(0);
      type_cast_2369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2369_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_116_2366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xix_xi28_2370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2376_inst_req_0;
      type_cast_2376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2376_inst_req_1;
      type_cast_2376_inst_ack_1<= rack(0);
      type_cast_2376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2376_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xix_xi28_2370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2376_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2399_inst_req_0;
      type_cast_2399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2399_inst_req_1;
      type_cast_2399_inst_ack_1<= rack(0);
      type_cast_2399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2399_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => torque_refx_x0_1920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xix_xi_2400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2506_inst_req_0;
      type_cast_2506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2506_inst_req_1;
      type_cast_2506_inst_ack_1<= rack(0);
      type_cast_2506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2506_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_153_2609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2506_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_82_2455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2512_inst_req_0;
      type_cast_2512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2512_inst_req_1;
      type_cast_2512_inst_ack_1<= rack(0);
      type_cast_2512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2512_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_152_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2512_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2540_inst_req_0;
      type_cast_2540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2540_inst_req_1;
      type_cast_2540_inst_ack_1<= rack(0);
      type_cast_2540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2540_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_183_2556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2540_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2542_inst_req_0;
      type_cast_2542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2542_inst_req_1;
      type_cast_2542_inst_ack_1<= rack(0);
      type_cast_2542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2542_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_85_2473,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2542_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2546_inst_req_0;
      type_cast_2546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2546_inst_req_1;
      type_cast_2546_inst_ack_1<= rack(0);
      type_cast_2546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2546_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_184_2562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2546_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2578_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2578_inst_req_0;
      type_cast_2578_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2578_inst_req_1;
      type_cast_2578_inst_ack_1<= rack(0);
      type_cast_2578_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2578_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_184_2562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2578_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2582_inst_req_0;
      type_cast_2582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2582_inst_req_1;
      type_cast_2582_inst_ack_1<= rack(0);
      type_cast_2582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2582_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_183_2556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2582_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2589_inst_req_0;
      type_cast_2589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2589_inst_req_1;
      type_cast_2589_inst_ack_1<= rack(0);
      type_cast_2589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2589_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_85_2473,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2589_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2591_inst_req_0;
      type_cast_2591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2591_inst_req_1;
      type_cast_2591_inst_ack_1<= rack(0);
      type_cast_2591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2591_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa7_2579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2591_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2598_inst_req_0;
      type_cast_2598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2598_inst_req_1;
      type_cast_2598_inst_ack_1<= rack(0);
      type_cast_2598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2598_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa8_2575,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2598_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2625_inst_req_0;
      type_cast_2625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2625_inst_req_1;
      type_cast_2625_inst_ack_1<= rack(0);
      type_cast_2625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2625_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_152_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2625_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2635_inst_req_0;
      type_cast_2635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2635_inst_req_1;
      type_cast_2635_inst_ack_1<= rack(0);
      type_cast_2635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2635_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa9_2622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2635_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2642_inst_req_0;
      type_cast_2642_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2642_inst_req_1;
      type_cast_2642_inst_ack_1<= rack(0);
      type_cast_2642_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2642_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_x0x_xix_xix_xi_2629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2642_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2644_inst_req_0;
      type_cast_2644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2644_inst_req_1;
      type_cast_2644_inst_ack_1<= rack(0);
      type_cast_2644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2644_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_82_2455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2644_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2683_inst_req_0;
      type_cast_2683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2683_inst_req_1;
      type_cast_2683_inst_ack_1<= rack(0);
      type_cast_2683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2683_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xix_xi_2730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2683_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2690_inst_req_0;
      type_cast_2690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2690_inst_req_1;
      type_cast_2690_inst_ack_1<= rack(0);
      type_cast_2690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2690_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_157_2699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2690_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2692_inst_req_0;
      type_cast_2692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2692_inst_req_1;
      type_cast_2692_inst_ack_1<= rack(0);
      type_cast_2692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2692_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi_2639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2692_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2741_inst_req_0;
      type_cast_2741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2741_inst_req_1;
      type_cast_2741_inst_ack_1<= rack(0);
      type_cast_2741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2741_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_157_2699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2741_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2745_inst_req_0;
      type_cast_2745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2745_inst_req_1;
      type_cast_2745_inst_ack_1<= rack(0);
      type_cast_2745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2745_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_156_2680,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2745_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2774_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2774_inst_req_0;
      type_cast_2774_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2774_inst_req_1;
      type_cast_2774_inst_ack_1<= rack(0);
      type_cast_2774_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2774_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xix_xi_2768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2774_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2776_inst_req_0;
      type_cast_2776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2776_inst_req_1;
      type_cast_2776_inst_ack_1<= rack(0);
      type_cast_2776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2776_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_88_2489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2776_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2780_inst_req_0;
      type_cast_2780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2780_inst_req_1;
      type_cast_2780_inst_ack_1<= rack(0);
      type_cast_2780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2780_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa6_2738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2780_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2782_inst_req_0;
      type_cast_2782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2782_inst_req_1;
      type_cast_2782_inst_ack_1<= rack(0);
      type_cast_2782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2782_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tempx_x0x_xphx_xix_xi_2639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2782_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2814_inst_req_0;
      type_cast_2814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2814_inst_req_1;
      type_cast_2814_inst_ack_1<= rack(0);
      type_cast_2814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2814_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_133_2811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xix_xi_2815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2821_inst_req_0;
      type_cast_2821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2821_inst_req_1;
      type_cast_2821_inst_ack_1<= rack(0);
      type_cast_2821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2821_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xix_xi_2815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2821_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2891_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2891_inst_req_0;
      type_cast_2891_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2891_inst_req_1;
      type_cast_2891_inst_ack_1<= rack(0);
      type_cast_2891_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2891_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_73_2859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2891_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2952_inst_req_0;
      type_cast_2952_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2952_inst_req_1;
      type_cast_2952_inst_ack_1<= rack(0);
      type_cast_2952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2952_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_97_2909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2952_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2962_inst_req_0;
      type_cast_2962_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2962_inst_req_1;
      type_cast_2962_inst_ack_1<= rack(0);
      type_cast_2962_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2962_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp10x_xi35x_xin_2949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10x_xi35_2963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2987_inst_req_0;
      type_cast_2987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2987_inst_req_1;
      type_cast_2987_inst_ack_1<= rack(0);
      type_cast_2987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2987_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_170_3093,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2987_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2989_inst_req_0;
      type_cast_2989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2989_inst_req_1;
      type_cast_2989_inst_ack_1<= rack(0);
      type_cast_2989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2989_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_120_2981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2989_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2993_inst_req_0;
      type_cast_2993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2993_inst_req_1;
      type_cast_2993_inst_ack_1<= rack(0);
      type_cast_2993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2993_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_169_3088,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3022_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3022_inst_req_0;
      type_cast_3022_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3022_inst_req_1;
      type_cast_3022_inst_ack_1<= rack(0);
      type_cast_3022_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3022_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_190_3039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3022_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3029_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3029_inst_req_0;
      type_cast_3029_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3029_inst_req_1;
      type_cast_3029_inst_ack_1<= rack(0);
      type_cast_3029_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3029_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_191_3045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3029_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3061_inst_req_0;
      type_cast_3061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3061_inst_req_1;
      type_cast_3061_inst_ack_1<= rack(0);
      type_cast_3061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3061_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_191_3045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3065_inst_req_0;
      type_cast_3065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3065_inst_req_1;
      type_cast_3065_inst_ack_1<= rack(0);
      type_cast_3065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3065_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_190_3039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3075_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3075_inst_req_0;
      type_cast_3075_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3075_inst_req_1;
      type_cast_3075_inst_ack_1<= rack(0);
      type_cast_3075_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3075_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa2_3062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3075_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3082_inst_req_0;
      type_cast_3082_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3082_inst_req_1;
      type_cast_3082_inst_ack_1<= rack(0);
      type_cast_3082_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3082_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa3_3058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3082_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3110_inst_req_0;
      type_cast_3110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3110_inst_req_1;
      type_cast_3110_inst_ack_1<= rack(0);
      type_cast_3110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3110_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_169_3088,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3110_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3173_inst_req_0;
      type_cast_3173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3173_inst_req_1;
      type_cast_3173_inst_ack_1<= rack(0);
      type_cast_3173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3173_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_3220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3173_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3180_inst_req_0;
      type_cast_3180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3180_inst_req_1;
      type_cast_3180_inst_ack_1<= rack(0);
      type_cast_3180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3180_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_212_3189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3180_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3182_inst_req_0;
      type_cast_3182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3182_inst_req_1;
      type_cast_3182_inst_ack_1<= rack(0);
      type_cast_3182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3182_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa4_3107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3182_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3231_inst_req_0;
      type_cast_3231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3231_inst_req_1;
      type_cast_3231_inst_ack_1<= rack(0);
      type_cast_3231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3231_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_212_3189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3231_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3235_inst_req_0;
      type_cast_3235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3235_inst_req_1;
      type_cast_3235_inst_ack_1<= rack(0);
      type_cast_3235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3235_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_211_3170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3235_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3253_inst_req_0;
      type_cast_3253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3253_inst_req_1;
      type_cast_3253_inst_ack_1<= rack(0);
      type_cast_3253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3253_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26x_xi_3247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3253_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3255_inst_req_0;
      type_cast_3255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3255_inst_req_1;
      type_cast_3255_inst_ack_1<= rack(0);
      type_cast_3255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3255_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_197_3135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3255_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3259_inst_req_0;
      type_cast_3259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3259_inst_req_1;
      type_cast_3259_inst_ack_1<= rack(0);
      type_cast_3259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3259_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa1_3228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3259_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3261_inst_req_0;
      type_cast_3261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3261_inst_req_1;
      type_cast_3261_inst_ack_1<= rack(0);
      type_cast_3261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3261_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa4_3107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3261_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3293_inst_req_0;
      type_cast_3293_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3293_inst_req_1;
      type_cast_3293_inst_ack_1<= rack(0);
      type_cast_3293_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3293_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_209_3290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3x_xi_3294,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3300_inst_req_0;
      type_cast_3300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3300_inst_req_1;
      type_cast_3300_inst_ack_1<= rack(0);
      type_cast_3300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3300_inst",
        buffer_size => 1,
        in_data_width => 32,
        out_data_width => 32
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3x_xi_3294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3300_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_1739_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_11_1738;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1739_branch_req_0,
          ack0 => if_stmt_1739_branch_ack_0,
          ack1 => if_stmt_1739_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1768_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_17_1767;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1768_branch_req_0,
          ack0 => if_stmt_1768_branch_ack_0,
          ack1 => if_stmt_1768_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1842_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_26_1841;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1842_branch_req_0,
          ack0 => if_stmt_1842_branch_ack_0,
          ack1 => if_stmt_1842_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1855_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_36_1854;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1855_branch_req_0,
          ack0 => if_stmt_1855_branch_ack_0,
          ack1 => if_stmt_1855_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1892_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_34_1891;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1892_branch_req_0,
          ack0 => if_stmt_1892_branch_ack_0,
          ack1 => if_stmt_1892_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1905_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_43_1904;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1905_branch_req_0,
          ack0 => if_stmt_1905_branch_ack_0,
          ack1 => if_stmt_1905_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1962_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_41_1961;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1962_branch_req_0,
          ack0 => if_stmt_1962_branch_ack_0,
          ack1 => if_stmt_1962_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2083_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_109_2082;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2083_branch_req_0,
          ack0 => if_stmt_2083_branch_ack_0,
          ack1 => if_stmt_2083_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2123_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_164_2122;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2123_branch_req_0,
          ack0 => if_stmt_2123_branch_ack_0,
          ack1 => if_stmt_2123_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2170_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_138_2169;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2170_branch_req_0,
          ack0 => if_stmt_2170_branch_ack_0,
          ack1 => if_stmt_2170_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2226_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xix_xi15_2225;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2226_branch_req_0,
          ack0 => if_stmt_2226_branch_ack_0,
          ack1 => if_stmt_2226_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2286_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xix_xi18_2279;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2286_branch_req_0,
          ack0 => if_stmt_2286_branch_ack_0,
          ack1 => if_stmt_2286_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2407_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_50_2406;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2407_branch_req_0,
          ack0 => if_stmt_2407_branch_ack_0,
          ack1 => if_stmt_2407_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2528_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_126_2527;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2528_branch_req_0,
          ack0 => if_stmt_2528_branch_ack_0,
          ack1 => if_stmt_2528_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2568_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_185_2567;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2568_branch_req_0,
          ack0 => if_stmt_2568_branch_ack_0,
          ack1 => if_stmt_2568_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2615_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_154_2614;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2615_branch_req_0,
          ack0 => if_stmt_2615_branch_ack_0,
          ack1 => if_stmt_2615_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2671_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xix_xi_2670;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2671_branch_req_0,
          ack0 => if_stmt_2671_branch_ack_0,
          ack1 => if_stmt_2671_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2731_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xix_xi_2724;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2731_branch_req_0,
          ack0 => if_stmt_2731_branch_ack_0,
          ack1 => if_stmt_2731_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2866_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_74_2865;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2866_branch_req_0,
          ack0 => if_stmt_2866_branch_ack_0,
          ack1 => if_stmt_2866_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2879_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_100_2878;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2879_branch_req_0,
          ack0 => if_stmt_2879_branch_ack_0,
          ack1 => if_stmt_2879_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2916_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_98_2915;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2916_branch_req_0,
          ack0 => if_stmt_2916_branch_ack_0,
          ack1 => if_stmt_2916_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2929_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_122_2928;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2929_branch_req_0,
          ack0 => if_stmt_2929_branch_ack_0,
          ack1 => if_stmt_2929_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2942_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_149_2941;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2942_branch_req_0,
          ack0 => if_stmt_2942_branch_ack_0,
          ack1 => if_stmt_2942_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3010_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_147_3009;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3010_branch_req_0,
          ack0 => if_stmt_3010_branch_ack_0,
          ack1 => if_stmt_3010_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3051_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_192_3050;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3051_branch_req_0,
          ack0 => if_stmt_3051_branch_ack_0,
          ack1 => if_stmt_3051_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3100_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_171_3099;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3100_branch_req_0,
          ack0 => if_stmt_3100_branch_ack_0,
          ack1 => if_stmt_3100_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3161_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond11x_xi_3160;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3161_branch_req_0,
          ack0 => if_stmt_3161_branch_ack_0,
          ack1 => if_stmt_3161_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3221_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xi_3214;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3221_branch_req_0,
          ack0 => if_stmt_3221_branch_ack_0,
          ack1 => if_stmt_3221_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2045_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2047_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2045_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_2045_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2045_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2050_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2045_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_2045_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2045_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_2047_wire_constant_cmp & expr_2050_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2045_branch_default_req_0,
          ack0 => switch_stmt_2045_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2490_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2492_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2490_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_2490_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2490_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_2495_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2490_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_2490_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_2490_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_2492_wire_constant_cmp & expr_2495_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_2490_branch_default_req_0,
          ack0 => switch_stmt_2490_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_f32_f32_1940_inst ADD_f32_f32_1830_inst ADD_f32_f32_1884_inst ADD_f32_f32_2835_inst ADD_f32_f32_2384_inst ADD_f32_f32_2395_inst ADD_f32_f32_1819_inst ADD_f32_f32_2908_inst ADD_f32_f32_2852_inst ADD_f32_f32_1809_inst 
    ApFloatAdd_group_0: Block -- 
      signal data_in: std_logic_vector(639 downto 0);
      signal data_out: std_logic_vector(319 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 9 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 9 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(9 downto 0) := (9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1, 4 => 1, 5 => 1, 6 => 1, 7 => 1, 8 => 1, 9 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_38_1936 & flux_rotor_prevx_x0_1690 & iNsTr_23_1826 & int_speed_err_prevx_x0_1704 & int_speed_errx_x0_1864 & iNsTr_32_1880 & iNsTr_68_2831 & flux_rotor_lpf_prevx_x0_1662 & iNsTr_46_2373 & iNsTr_10_1733 & iNsTr_48_2391 & theta_prevx_x0_1683 & iNsTr_21_1815 & speed_err_prevx_x0_1676 & int_flux_errx_x0_2888 & iNsTr_96_2904 & iNsTr_71_2848 & int_flux_err_temp_2x_x0_1669 & iNsTr_19_1805 & spd_lpf_prevx_x0_1697;
      iNsTr_39_1941 <= data_out(319 downto 288);
      iNsTr_24_1831 <= data_out(287 downto 256);
      iNsTr_33_1885 <= data_out(255 downto 224);
      iNsTr_69_2836 <= data_out(223 downto 192);
      iNsTr_47_2385 <= data_out(191 downto 160);
      iNsTr_49_2396 <= data_out(159 downto 128);
      iNsTr_22_1820 <= data_out(127 downto 96);
      iNsTr_97_2909 <= data_out(95 downto 64);
      iNsTr_72_2853 <= data_out(63 downto 32);
      iNsTr_20_1810 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      reqL_unguarded(9) <= ADD_f32_f32_1940_inst_req_0;
      reqL_unguarded(8) <= ADD_f32_f32_1830_inst_req_0;
      reqL_unguarded(7) <= ADD_f32_f32_1884_inst_req_0;
      reqL_unguarded(6) <= ADD_f32_f32_2835_inst_req_0;
      reqL_unguarded(5) <= ADD_f32_f32_2384_inst_req_0;
      reqL_unguarded(4) <= ADD_f32_f32_2395_inst_req_0;
      reqL_unguarded(3) <= ADD_f32_f32_1819_inst_req_0;
      reqL_unguarded(2) <= ADD_f32_f32_2908_inst_req_0;
      reqL_unguarded(1) <= ADD_f32_f32_2852_inst_req_0;
      reqL_unguarded(0) <= ADD_f32_f32_1809_inst_req_0;
      ADD_f32_f32_1940_inst_ack_0 <= ackL_unguarded(9);
      ADD_f32_f32_1830_inst_ack_0 <= ackL_unguarded(8);
      ADD_f32_f32_1884_inst_ack_0 <= ackL_unguarded(7);
      ADD_f32_f32_2835_inst_ack_0 <= ackL_unguarded(6);
      ADD_f32_f32_2384_inst_ack_0 <= ackL_unguarded(5);
      ADD_f32_f32_2395_inst_ack_0 <= ackL_unguarded(4);
      ADD_f32_f32_1819_inst_ack_0 <= ackL_unguarded(3);
      ADD_f32_f32_2908_inst_ack_0 <= ackL_unguarded(2);
      ADD_f32_f32_2852_inst_ack_0 <= ackL_unguarded(1);
      ADD_f32_f32_1809_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(9) <= ADD_f32_f32_1940_inst_req_1;
      reqR_unguarded(8) <= ADD_f32_f32_1830_inst_req_1;
      reqR_unguarded(7) <= ADD_f32_f32_1884_inst_req_1;
      reqR_unguarded(6) <= ADD_f32_f32_2835_inst_req_1;
      reqR_unguarded(5) <= ADD_f32_f32_2384_inst_req_1;
      reqR_unguarded(4) <= ADD_f32_f32_2395_inst_req_1;
      reqR_unguarded(3) <= ADD_f32_f32_1819_inst_req_1;
      reqR_unguarded(2) <= ADD_f32_f32_2908_inst_req_1;
      reqR_unguarded(1) <= ADD_f32_f32_2852_inst_req_1;
      reqR_unguarded(0) <= ADD_f32_f32_1809_inst_req_1;
      ADD_f32_f32_1940_inst_ack_1 <= ackR_unguarded(9);
      ADD_f32_f32_1830_inst_ack_1 <= ackR_unguarded(8);
      ADD_f32_f32_1884_inst_ack_1 <= ackR_unguarded(7);
      ADD_f32_f32_2835_inst_ack_1 <= ackR_unguarded(6);
      ADD_f32_f32_2384_inst_ack_1 <= ackR_unguarded(5);
      ADD_f32_f32_2395_inst_ack_1 <= ackR_unguarded(4);
      ADD_f32_f32_1819_inst_ack_1 <= ackR_unguarded(3);
      ADD_f32_f32_2908_inst_ack_1 <= ackR_unguarded(2);
      ADD_f32_f32_2852_inst_ack_1 <= ackR_unguarded(1);
      ADD_f32_f32_1809_inst_ack_1 <= ackR_unguarded(0);
      ApFloatAdd_group_0_accessRegulator_0: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_1: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_2: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_3: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_4: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_5: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_6: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_7: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_8: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_0_accessRegulator_9: access_regulator_base generic map (name => "ApFloatAdd_group_0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 10, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatAdd_group_0",
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 10,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_f64_f64_1755_inst ADD_f64_f64_1783_inst 
    ApFloatAdd_group_1: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 1, 1 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_13_1750 & type_cast_1754_wire_constant & iNsTr_28_1778 & type_cast_1782_wire_constant;
      iNsTr_14_1756 <= data_out(127 downto 64);
      iNsTr_29_1784 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      reqL_unguarded(1) <= ADD_f64_f64_1755_inst_req_0;
      reqL_unguarded(0) <= ADD_f64_f64_1783_inst_req_0;
      ADD_f64_f64_1755_inst_ack_0 <= ackL_unguarded(1);
      ADD_f64_f64_1783_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ADD_f64_f64_1755_inst_req_1;
      reqR_unguarded(0) <= ADD_f64_f64_1783_inst_req_1;
      ADD_f64_f64_1755_inst_ack_1 <= ackR_unguarded(1);
      ADD_f64_f64_1783_inst_ack_1 <= ackR_unguarded(0);
      ApFloatAdd_group_1_accessRegulator_0: access_regulator_base generic map (name => "ApFloatAdd_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatAdd_group_1_accessRegulator_1: access_regulator_base generic map (name => "ApFloatAdd_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 2, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatAdd_group_1",
          operator_id => "ApFloatAdd",
          exponent_width => 11,
          fraction_width => 52, 
          no_arbitration => false,
          num_reqs => 2,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u32_u32_2158_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xix_xi10_2147 & quotientx_x05x_xix_xix_xi4_2064;
      iNsTr_136_2159 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2158_inst_req_0;
      ADD_u32_u32_2158_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2158_inst_req_1;
      ADD_u32_u32_2158_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u32_u32_2284_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_140_2235;
      indvarx_xnextx_xix_xi19_2285 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2284_inst_req_0;
      ADD_u32_u32_2284_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2284_inst_req_1;
      ADD_u32_u32_2284_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ADD_u32_u32_2317_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp21x_xix_xi22_2313 & iNsTr_53_1980;
      tmp25x_xix_xi23_2318 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2317_inst_req_0;
      ADD_u32_u32_2317_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2317_inst_req_1;
      ADD_u32_u32_2317_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ADD_u32_u32_2355_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_113_2350;
      iNsTr_114_2356 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2355_inst_req_0;
      ADD_u32_u32_2355_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2355_inst_req_1;
      ADD_u32_u32_2355_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : ADD_u32_u32_2603_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xix_xi_2592 & quotientx_x05x_xix_xix_xi_2509;
      iNsTr_152_2604 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2603_inst_req_0;
      ADD_u32_u32_2603_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2603_inst_req_1;
      ADD_u32_u32_2603_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ADD_u32_u32_2729_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_156_2680;
      indvarx_xnextx_xix_xi_2730 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2729_inst_req_0;
      ADD_u32_u32_2729_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2729_inst_req_1;
      ADD_u32_u32_2729_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ADD_u32_u32_2762_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_77_2425 & tmp21x_xix_xi_2758;
      tmp25x_xix_xi_2763 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2762_inst_req_0;
      ADD_u32_u32_2762_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2762_inst_req_1;
      ADD_u32_u32_2762_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ADD_u32_u32_2800_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_130_2795;
      iNsTr_131_2801 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2800_inst_req_0;
      ADD_u32_u32_2800_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2800_inst_req_1;
      ADD_u32_u32_2800_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ADD_u32_u32_3087_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x0x_xlcssax_xix_xi_3076 & quotientx_x05x_xix_xi_2990;
      iNsTr_169_3088 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3087_inst_req_0;
      ADD_u32_u32_3087_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3087_inst_req_1;
      ADD_u32_u32_3087_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ADD_u32_u32_3134_inst 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_196_3129;
      iNsTr_197_3135 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3134_inst_req_0;
      ADD_u32_u32_3134_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3134_inst_req_1;
      ADD_u32_u32_3134_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111110000010",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ADD_u32_u32_3219_inst 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_211_3170;
      indvarx_xnextx_xi_3220 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3219_inst_req_0;
      ADD_u32_u32_3219_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3219_inst_req_1;
      ADD_u32_u32_3219_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ADD_u32_u32_3241_inst 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_196_3129;
      tmp25x_xi_3242 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3241_inst_req_0;
      ADD_u32_u32_3241_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3241_inst_req_1;
      ADD_u32_u32_3241_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111110000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ADD_u32_u32_3279_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_206_3274;
      iNsTr_207_3280 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_3279_inst_req_0;
      ADD_u32_u32_3279_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_3279_inst_req_1;
      ADD_u32_u32_3279_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000100000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : AND_u1_u1_2224_inst 
    ApIntAnd_group_15: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_93_2212 & iNsTr_94_2220;
      orx_xcond11x_xix_xi15_2225 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2224_inst_req_0;
      AND_u1_u1_2224_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2224_inst_req_1;
      AND_u1_u1_2224_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : AND_u1_u1_2278_inst 
    ApIntAnd_group_16: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_143_2266 & iNsTr_144_2274;
      orx_xcondx_xix_xi18_2279 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2278_inst_req_0;
      AND_u1_u1_2278_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2278_inst_req_1;
      AND_u1_u1_2278_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : AND_u1_u1_2669_inst 
    ApIntAnd_group_17: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_105_2657 & iNsTr_106_2665;
      orx_xcond11x_xix_xi_2670 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2669_inst_req_0;
      AND_u1_u1_2669_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2669_inst_req_1;
      AND_u1_u1_2669_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : AND_u1_u1_2723_inst 
    ApIntAnd_group_18: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_159_2711 & iNsTr_160_2719;
      orx_xcondx_xix_xi_2724 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2723_inst_req_0;
      AND_u1_u1_2723_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2723_inst_req_1;
      AND_u1_u1_2723_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : AND_u1_u1_3159_inst 
    ApIntAnd_group_19: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_199_3147 & iNsTr_200_3155;
      orx_xcond11x_xi_3160 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3159_inst_req_0;
      AND_u1_u1_3159_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3159_inst_req_1;
      AND_u1_u1_3159_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : AND_u1_u1_3213_inst 
    ApIntAnd_group_20: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_214_3201 & iNsTr_215_3209;
      orx_xcondx_xi_3214 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3213_inst_req_0;
      AND_u1_u1_3213_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3213_inst_req_1;
      AND_u1_u1_3213_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : AND_u32_u32_1979_inst 
    ApIntAnd_group_21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_52_1974;
      iNsTr_53_1980 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_1979_inst_req_0;
      AND_u32_u32_1979_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_1979_inst_req_1;
      AND_u32_u32_1979_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : AND_u32_u32_1991_inst 
    ApIntAnd_group_22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_54_1986;
      iNsTr_55_1992 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_1991_inst_req_0;
      AND_u32_u32_1991_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_1991_inst_req_1;
      AND_u32_u32_1991_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : AND_u32_u32_2003_inst 
    ApIntAnd_group_23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_56_1998;
      iNsTr_57_2004 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2003_inst_req_0;
      AND_u32_u32_2003_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2003_inst_req_1;
      AND_u32_u32_2003_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : AND_u32_u32_2021_inst 
    ApIntAnd_group_24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_59_2016;
      iNsTr_60_2022 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2021_inst_req_0;
      AND_u32_u32_2021_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2021_inst_req_1;
      AND_u32_u32_2021_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : AND_u32_u32_2038_inst 
    ApIntAnd_group_25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_62_2033;
      iNsTr_63_2039 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2038_inst_req_0;
      AND_u32_u32_2038_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2038_inst_req_1;
      AND_u32_u32_2038_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : AND_u32_u32_2205_inst 
    ApIntAnd_group_26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi14_2194;
      iNsTr_92_2206 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2205_inst_req_0;
      AND_u32_u32_2205_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2205_inst_req_1;
      AND_u32_u32_2205_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : AND_u32_u32_2259_inst 
    ApIntAnd_group_27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_141_2254;
      iNsTr_142_2260 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2259_inst_req_0;
      AND_u32_u32_2259_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2259_inst_req_1;
      AND_u32_u32_2259_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : AND_u32_u32_2343_inst 
    ApIntAnd_group_28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xix_xi27_2332;
      iNsTr_112_2344 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2343_inst_req_0;
      AND_u32_u32_2343_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2343_inst_req_1;
      AND_u32_u32_2343_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : AND_u32_u32_2424_inst 
    ApIntAnd_group_29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_76_2419;
      iNsTr_77_2425 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2424_inst_req_0;
      AND_u32_u32_2424_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2424_inst_req_1;
      AND_u32_u32_2424_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : AND_u32_u32_2436_inst 
    ApIntAnd_group_30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_78_2431;
      iNsTr_79_2437 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2436_inst_req_0;
      AND_u32_u32_2436_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2436_inst_req_1;
      AND_u32_u32_2436_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : AND_u32_u32_2448_inst 
    ApIntAnd_group_31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_80_2443;
      iNsTr_81_2449 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2448_inst_req_0;
      AND_u32_u32_2448_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2448_inst_req_1;
      AND_u32_u32_2448_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : AND_u32_u32_2466_inst 
    ApIntAnd_group_32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_83_2461;
      iNsTr_84_2467 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2466_inst_req_0;
      AND_u32_u32_2466_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2466_inst_req_1;
      AND_u32_u32_2466_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : AND_u32_u32_2483_inst 
    ApIntAnd_group_33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_86_2478;
      iNsTr_87_2484 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2483_inst_req_0;
      AND_u32_u32_2483_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2483_inst_req_1;
      AND_u32_u32_2483_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : AND_u32_u32_2650_inst 
    ApIntAnd_group_34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi_2639;
      iNsTr_104_2651 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2650_inst_req_0;
      AND_u32_u32_2650_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2650_inst_req_1;
      AND_u32_u32_2650_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : AND_u32_u32_2704_inst 
    ApIntAnd_group_35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_157_2699;
      iNsTr_158_2705 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2704_inst_req_0;
      AND_u32_u32_2704_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2704_inst_req_1;
      AND_u32_u32_2704_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : AND_u32_u32_2788_inst 
    ApIntAnd_group_36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xix_xi_2777;
      iNsTr_129_2789 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2788_inst_req_0;
      AND_u32_u32_2788_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2788_inst_req_1;
      AND_u32_u32_2788_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : AND_u32_u32_2974_inst 
    ApIntAnd_group_37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_118_2969;
      iNsTr_119_2975 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_2974_inst_req_0;
      AND_u32_u32_2974_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_2974_inst_req_1;
      AND_u32_u32_2974_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00111111111111111111111110000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : AND_u32_u32_3122_inst 
    ApIntAnd_group_38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi35_2963;
      iNsTr_195_3123 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3122_inst_req_0;
      AND_u32_u32_3122_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3122_inst_req_1;
      AND_u32_u32_3122_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "10000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : AND_u32_u32_3128_inst 
    ApIntAnd_group_39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_194_3117;
      iNsTr_196_3129 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3128_inst_req_0;
      AND_u32_u32_3128_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3128_inst_req_1;
      AND_u32_u32_3128_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : AND_u32_u32_3140_inst 
    ApIntAnd_group_40: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa4_3107;
      iNsTr_198_3141 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3140_inst_req_0;
      AND_u32_u32_3140_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3140_inst_req_1;
      AND_u32_u32_3140_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : AND_u32_u32_3194_inst 
    ApIntAnd_group_41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_212_3189;
      iNsTr_213_3195 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3194_inst_req_0;
      AND_u32_u32_3194_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3194_inst_req_1;
      AND_u32_u32_3194_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : AND_u32_u32_3267_inst 
    ApIntAnd_group_42: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xlcssax_xi_3256;
      iNsTr_205_3268 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_3267_inst_req_0;
      AND_u32_u32_3267_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_3267_inst_req_1;
      AND_u32_u32_3267_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000011111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : EQ_f32_u1_1960_inst 
    ApFloatUeq_group_43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_40_1947;
      iNsTr_41_1961 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_1960_inst_req_0;
      EQ_f32_u1_1960_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_1960_inst_req_1;
      EQ_f32_u1_1960_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_43",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : EQ_f32_u1_2405_inst 
    ApFloatUeq_group_44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= torque_refx_x0_1920;
      iNsTr_50_2406 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_2405_inst_req_0;
      EQ_f32_u1_2405_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_2405_inst_req_1;
      EQ_f32_u1_2405_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_44",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : EQ_f32_u1_2940_inst 
    ApFloatUeq_group_45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_97_2909;
      iNsTr_149_2941 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_f32_u1_2940_inst_req_0;
      EQ_f32_u1_2940_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_f32_u1_2940_inst_req_1;
      EQ_f32_u1_2940_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUeq",
          name => "ApFloatUeq_group_45",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : EQ_u32_u1_2211_inst 
    ApIntEq_group_46: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_92_2206;
      iNsTr_93_2212 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2211_inst_req_0;
      EQ_u32_u1_2211_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2211_inst_req_1;
      EQ_u32_u1_2211_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : EQ_u32_u1_2265_inst 
    ApIntEq_group_47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_142_2260;
      iNsTr_143_2266 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2265_inst_req_0;
      EQ_u32_u1_2265_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2265_inst_req_1;
      EQ_u32_u1_2265_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : EQ_u32_u1_2656_inst 
    ApIntEq_group_48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_104_2651;
      iNsTr_105_2657 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2656_inst_req_0;
      EQ_u32_u1_2656_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2656_inst_req_1;
      EQ_u32_u1_2656_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : EQ_u32_u1_2710_inst 
    ApIntEq_group_49: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_158_2705;
      iNsTr_159_2711 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2710_inst_req_0;
      EQ_u32_u1_2710_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2710_inst_req_1;
      EQ_u32_u1_2710_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : EQ_u32_u1_3146_inst 
    ApIntEq_group_50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_198_3141;
      iNsTr_199_3147 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3146_inst_req_0;
      EQ_u32_u1_3146_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3146_inst_req_1;
      EQ_u32_u1_3146_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : EQ_u32_u1_3200_inst 
    ApIntEq_group_51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_213_3195;
      iNsTr_214_3201 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_3200_inst_req_0;
      EQ_u32_u1_3200_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_3200_inst_req_1;
      EQ_u32_u1_3200_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : LSHR_u32_u32_1973_inst 
    ApIntLSHR_group_52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi1_1951;
      iNsTr_52_1974 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_1973_inst_req_0;
      LSHR_u32_u32_1973_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_1973_inst_req_1;
      LSHR_u32_u32_1973_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : LSHR_u32_u32_1985_inst 
    ApIntLSHR_group_53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_1955;
      iNsTr_54_1986 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_1985_inst_req_0;
      LSHR_u32_u32_1985_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_1985_inst_req_1;
      LSHR_u32_u32_1985_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : LSHR_u32_u32_2015_inst 
    ApIntLSHR_group_54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_1955;
      iNsTr_59_2016 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2015_inst_req_0;
      LSHR_u32_u32_2015_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2015_inst_req_1;
      LSHR_u32_u32_2015_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : LSHR_u32_u32_2076_inst 
    ApIntLSHR_group_55: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi3_2058;
      iNsTr_108_2077 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2076_inst_req_0;
      LSHR_u32_u32_2076_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2076_inst_req_1;
      LSHR_u32_u32_2076_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_55",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : LSHR_u32_u32_2418_inst 
    ApIntLSHR_group_56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi_2400;
      iNsTr_76_2419 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2418_inst_req_0;
      LSHR_u32_u32_2418_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2418_inst_req_1;
      LSHR_u32_u32_2418_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_56",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : LSHR_u32_u32_2430_inst 
    ApIntLSHR_group_57: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_1955;
      iNsTr_78_2431 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2430_inst_req_0;
      LSHR_u32_u32_2430_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2430_inst_req_1;
      LSHR_u32_u32_2430_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : LSHR_u32_u32_2460_inst 
    ApIntLSHR_group_58: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_1955;
      iNsTr_83_2461 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2460_inst_req_0;
      LSHR_u32_u32_2460_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2460_inst_req_1;
      LSHR_u32_u32_2460_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : LSHR_u32_u32_2521_inst 
    ApIntLSHR_group_59: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi_2503;
      iNsTr_125_2522 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_2521_inst_req_0;
      LSHR_u32_u32_2521_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_2521_inst_req_1;
      LSHR_u32_u32_2521_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : LSHR_u32_u32_3002_inst 
    ApIntLSHR_group_60: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xi_2984;
      iNsTr_146_3003 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3002_inst_req_0;
      LSHR_u32_u32_3002_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3002_inst_req_1;
      LSHR_u32_u32_3002_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : LSHR_u32_u32_3116_inst 
    ApIntLSHR_group_61: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi35_2963;
      iNsTr_194_3117 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_3116_inst_req_0;
      LSHR_u32_u32_3116_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_3116_inst_req_1;
      LSHR_u32_u32_3116_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : MUL_f32_f32_1916_inst MUL_f32_f32_1935_inst MUL_f32_f32_1825_inst MUL_f32_f32_1879_inst MUL_f32_f32_1946_inst MUL_f32_f32_2390_inst MUL_f32_f32_2858_inst MUL_f32_f32_2830_inst MUL_f32_f32_2903_inst MUL_f32_f32_2847_inst MUL_f32_f32_1804_inst MUL_f32_f32_3321_inst MUL_f32_f32_3327_inst MUL_f32_f32_3333_inst 
    ApFloatMul_group_62: Block -- 
      signal data_in: std_logic_vector(895 downto 0);
      signal data_out: std_logic_vector(447 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1, 4 => 1, 5 => 1, 6 => 1, 7 => 1, 8 => 1, 9 => 1, 10 => 1, 11 => 1, 12 => 1, 13 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_33_1885 & type_cast_1915_wire_constant & iNsTr_2_1721 & type_cast_1934_wire_constant & iNsTr_22_1820 & type_cast_1824_wire_constant & iNsTr_21_1815 & type_cast_1878_wire_constant & iNsTr_4_1724 & type_cast_1945_wire_constant & iNsTr_47_2385 & type_cast_2389_wire_constant & iNsTr_72_2853 & type_cast_2857_wire_constant & iNsTr_39_1941 & type_cast_2829_wire_constant & iNsTr_70_2842 & type_cast_2902_wire_constant & iNsTr_70_2842 & type_cast_2846_wire_constant & iNsTr_6_1727 & type_cast_1803_wire_constant & iNsTr_20_1810 & type_cast_3320_wire_constant & iNsTr_39_1941 & type_cast_3326_wire_constant & iNsTr_69_2836 & type_cast_3332_wire_constant;
      phitmp32_1917 <= data_out(447 downto 416);
      iNsTr_38_1936 <= data_out(415 downto 384);
      iNsTr_23_1826 <= data_out(383 downto 352);
      iNsTr_32_1880 <= data_out(351 downto 320);
      iNsTr_40_1947 <= data_out(319 downto 288);
      iNsTr_48_2391 <= data_out(287 downto 256);
      iNsTr_73_2859 <= data_out(255 downto 224);
      iNsTr_68_2831 <= data_out(223 downto 192);
      iNsTr_96_2904 <= data_out(191 downto 160);
      iNsTr_71_2848 <= data_out(159 downto 128);
      iNsTr_19_1805 <= data_out(127 downto 96);
      phitmp_3322 <= data_out(95 downto 64);
      phitmp31_3328 <= data_out(63 downto 32);
      phitmp33_3334 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      reqL_unguarded(13) <= MUL_f32_f32_1916_inst_req_0;
      reqL_unguarded(12) <= MUL_f32_f32_1935_inst_req_0;
      reqL_unguarded(11) <= MUL_f32_f32_1825_inst_req_0;
      reqL_unguarded(10) <= MUL_f32_f32_1879_inst_req_0;
      reqL_unguarded(9) <= MUL_f32_f32_1946_inst_req_0;
      reqL_unguarded(8) <= MUL_f32_f32_2390_inst_req_0;
      reqL_unguarded(7) <= MUL_f32_f32_2858_inst_req_0;
      reqL_unguarded(6) <= MUL_f32_f32_2830_inst_req_0;
      reqL_unguarded(5) <= MUL_f32_f32_2903_inst_req_0;
      reqL_unguarded(4) <= MUL_f32_f32_2847_inst_req_0;
      reqL_unguarded(3) <= MUL_f32_f32_1804_inst_req_0;
      reqL_unguarded(2) <= MUL_f32_f32_3321_inst_req_0;
      reqL_unguarded(1) <= MUL_f32_f32_3327_inst_req_0;
      reqL_unguarded(0) <= MUL_f32_f32_3333_inst_req_0;
      MUL_f32_f32_1916_inst_ack_0 <= ackL_unguarded(13);
      MUL_f32_f32_1935_inst_ack_0 <= ackL_unguarded(12);
      MUL_f32_f32_1825_inst_ack_0 <= ackL_unguarded(11);
      MUL_f32_f32_1879_inst_ack_0 <= ackL_unguarded(10);
      MUL_f32_f32_1946_inst_ack_0 <= ackL_unguarded(9);
      MUL_f32_f32_2390_inst_ack_0 <= ackL_unguarded(8);
      MUL_f32_f32_2858_inst_ack_0 <= ackL_unguarded(7);
      MUL_f32_f32_2830_inst_ack_0 <= ackL_unguarded(6);
      MUL_f32_f32_2903_inst_ack_0 <= ackL_unguarded(5);
      MUL_f32_f32_2847_inst_ack_0 <= ackL_unguarded(4);
      MUL_f32_f32_1804_inst_ack_0 <= ackL_unguarded(3);
      MUL_f32_f32_3321_inst_ack_0 <= ackL_unguarded(2);
      MUL_f32_f32_3327_inst_ack_0 <= ackL_unguarded(1);
      MUL_f32_f32_3333_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= MUL_f32_f32_1916_inst_req_1;
      reqR_unguarded(12) <= MUL_f32_f32_1935_inst_req_1;
      reqR_unguarded(11) <= MUL_f32_f32_1825_inst_req_1;
      reqR_unguarded(10) <= MUL_f32_f32_1879_inst_req_1;
      reqR_unguarded(9) <= MUL_f32_f32_1946_inst_req_1;
      reqR_unguarded(8) <= MUL_f32_f32_2390_inst_req_1;
      reqR_unguarded(7) <= MUL_f32_f32_2858_inst_req_1;
      reqR_unguarded(6) <= MUL_f32_f32_2830_inst_req_1;
      reqR_unguarded(5) <= MUL_f32_f32_2903_inst_req_1;
      reqR_unguarded(4) <= MUL_f32_f32_2847_inst_req_1;
      reqR_unguarded(3) <= MUL_f32_f32_1804_inst_req_1;
      reqR_unguarded(2) <= MUL_f32_f32_3321_inst_req_1;
      reqR_unguarded(1) <= MUL_f32_f32_3327_inst_req_1;
      reqR_unguarded(0) <= MUL_f32_f32_3333_inst_req_1;
      MUL_f32_f32_1916_inst_ack_1 <= ackR_unguarded(13);
      MUL_f32_f32_1935_inst_ack_1 <= ackR_unguarded(12);
      MUL_f32_f32_1825_inst_ack_1 <= ackR_unguarded(11);
      MUL_f32_f32_1879_inst_ack_1 <= ackR_unguarded(10);
      MUL_f32_f32_1946_inst_ack_1 <= ackR_unguarded(9);
      MUL_f32_f32_2390_inst_ack_1 <= ackR_unguarded(8);
      MUL_f32_f32_2858_inst_ack_1 <= ackR_unguarded(7);
      MUL_f32_f32_2830_inst_ack_1 <= ackR_unguarded(6);
      MUL_f32_f32_2903_inst_ack_1 <= ackR_unguarded(5);
      MUL_f32_f32_2847_inst_ack_1 <= ackR_unguarded(4);
      MUL_f32_f32_1804_inst_ack_1 <= ackR_unguarded(3);
      MUL_f32_f32_3321_inst_ack_1 <= ackR_unguarded(2);
      MUL_f32_f32_3327_inst_ack_1 <= ackR_unguarded(1);
      MUL_f32_f32_3333_inst_ack_1 <= ackR_unguarded(0);
      ApFloatMul_group_62_accessRegulator_0: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_1: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_2: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_3: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_4: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_5: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_6: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_7: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_8: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_9: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_10: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_11: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_12: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_62_accessRegulator_13: access_regulator_base generic map (name => "ApFloatMul_group_62_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 14, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatMul_group_62",
          operator_id => "ApFloatMul",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 14,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : NEQ_i32_u1_2219_inst 
    ApIntNe_group_63: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2215_wire;
      iNsTr_94_2220 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2219_inst_req_0;
      NEQ_i32_u1_2219_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2219_inst_req_1;
      NEQ_i32_u1_2219_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : NEQ_i32_u1_2273_inst 
    ApIntNe_group_64: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2269_wire;
      iNsTr_144_2274 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2273_inst_req_0;
      NEQ_i32_u1_2273_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2273_inst_req_1;
      NEQ_i32_u1_2273_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : NEQ_i32_u1_2664_inst 
    ApIntNe_group_65: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2660_wire;
      iNsTr_106_2665 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2664_inst_req_0;
      NEQ_i32_u1_2664_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2664_inst_req_1;
      NEQ_i32_u1_2664_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : NEQ_i32_u1_2718_inst 
    ApIntNe_group_66: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2714_wire;
      iNsTr_160_2719 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_2718_inst_req_0;
      NEQ_i32_u1_2718_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_2718_inst_req_1;
      NEQ_i32_u1_2718_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : NEQ_i32_u1_3154_inst 
    ApIntNe_group_67: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3150_wire;
      iNsTr_200_3155 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3154_inst_req_0;
      NEQ_i32_u1_3154_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3154_inst_req_1;
      NEQ_i32_u1_3154_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : NEQ_i32_u1_3208_inst 
    ApIntNe_group_68: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= type_cast_3204_wire;
      iNsTr_215_3209 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NEQ_i32_u1_3208_inst_req_0;
      NEQ_i32_u1_3208_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NEQ_i32_u1_3208_inst_req_1;
      NEQ_i32_u1_3208_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          name => "ApIntNe_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : OR_u32_u32_2009_inst 
    ApIntOr_group_69: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_57_2004;
      iNsTr_58_2010 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2009_inst_req_0;
      OR_u32_u32_2009_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2009_inst_req_1;
      OR_u32_u32_2009_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : OR_u32_u32_2027_inst 
    ApIntOr_group_70: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_60_2022;
      iNsTr_61_2028 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2027_inst_req_0;
      OR_u32_u32_2027_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2027_inst_req_1;
      OR_u32_u32_2027_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000010000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : OR_u32_u32_2306_inst 
    ApIntOr_group_71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_54_1986;
      xx_xnotx_xi21_2307 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2306_inst_req_0;
      OR_u32_u32_2306_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2306_inst_req_1;
      OR_u32_u32_2306_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111100000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : OR_u32_u32_2360_inst 
    ApIntOr_group_72: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_112_2344 & iNsTr_63_2039;
      iNsTr_115_2361 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2360_inst_req_0;
      OR_u32_u32_2360_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2360_inst_req_1;
      OR_u32_u32_2360_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : OR_u32_u32_2365_inst 
    ApIntOr_group_73: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_115_2361 & iNsTr_114_2356;
      iNsTr_116_2366 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2365_inst_req_0;
      OR_u32_u32_2365_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2365_inst_req_1;
      OR_u32_u32_2365_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : OR_u32_u32_2454_inst 
    ApIntOr_group_74: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_81_2449;
      iNsTr_82_2455 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2454_inst_req_0;
      OR_u32_u32_2454_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2454_inst_req_1;
      OR_u32_u32_2454_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_74",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : OR_u32_u32_2472_inst 
    ApIntOr_group_75: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_84_2467;
      iNsTr_85_2473 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2472_inst_req_0;
      OR_u32_u32_2472_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2472_inst_req_1;
      OR_u32_u32_2472_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_75",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000010000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : OR_u32_u32_2751_inst 
    ApIntOr_group_76: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_78_2431;
      xx_xnotx_xi_2752 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2751_inst_req_0;
      OR_u32_u32_2751_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2751_inst_req_1;
      OR_u32_u32_2751_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_76",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111100000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : OR_u32_u32_2805_inst 
    ApIntOr_group_77: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_129_2789 & iNsTr_87_2484;
      iNsTr_132_2806 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2805_inst_req_0;
      OR_u32_u32_2805_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2805_inst_req_1;
      OR_u32_u32_2805_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_77",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : OR_u32_u32_2810_inst 
    ApIntOr_group_78: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_132_2806 & iNsTr_131_2801;
      iNsTr_133_2811 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2810_inst_req_0;
      OR_u32_u32_2810_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2810_inst_req_1;
      OR_u32_u32_2810_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_78",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : OR_u32_u32_2980_inst 
    ApIntOr_group_79: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_119_2975;
      iNsTr_120_2981 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_2980_inst_req_0;
      OR_u32_u32_2980_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_2980_inst_req_1;
      OR_u32_u32_2980_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_79",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : OR_u32_u32_3284_inst 
    ApIntOr_group_80: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_207_3280 & iNsTr_195_3123;
      iNsTr_208_3285 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3284_inst_req_0;
      OR_u32_u32_3284_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3284_inst_req_1;
      OR_u32_u32_3284_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_80",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : OR_u32_u32_3289_inst 
    ApIntOr_group_81: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_208_3285 & iNsTr_205_3268;
      iNsTr_209_3290 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_3289_inst_req_0;
      OR_u32_u32_3289_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_3289_inst_req_1;
      OR_u32_u32_3289_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_81",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : SGT_f32_u1_1766_inst 
    ApFloatUgt_group_82: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= speed_refx_x1_1711 & iNsTr_8_1730;
      iNsTr_17_1767 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_1766_inst_req_0;
      SGT_f32_u1_1766_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_1766_inst_req_1;
      SGT_f32_u1_1766_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_82",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : SGT_f32_u1_1903_inst 
    ApFloatUgt_group_83: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_33_1885;
      iNsTr_43_1904 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_1903_inst_req_0;
      SGT_f32_u1_1903_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_1903_inst_req_1;
      SGT_f32_u1_1903_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_83",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01000001101000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : SGT_f32_u1_2877_inst 
    ApFloatUgt_group_84: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_73_2859;
      iNsTr_100_2878 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_2877_inst_req_0;
      SGT_f32_u1_2877_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_2877_inst_req_1;
      SGT_f32_u1_2877_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_84",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00111111100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : SGT_f32_u1_2927_inst 
    ApFloatUgt_group_85: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_97_2909;
      iNsTr_122_2928 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f32_u1_2927_inst_req_0;
      SGT_f32_u1_2927_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f32_u1_2927_inst_req_1;
      SGT_f32_u1_2927_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_85",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : SGT_f64_u1_1853_inst 
    ApFloatUgt_group_86: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_25_1835;
      iNsTr_36_1854 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_1853_inst_req_0;
      SGT_f64_u1_1853_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_1853_inst_req_1;
      SGT_f64_u1_1853_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_86",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0100000000100100000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : SHL_u32_u32_1997_inst 
    ApIntSHL_group_87: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi1_1951;
      iNsTr_56_1998 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_1997_inst_req_0;
      SHL_u32_u32_1997_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_1997_inst_req_1;
      SHL_u32_u32_1997_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_87",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : SHL_u32_u32_2110_inst 
    ApIntSHL_group_88: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xix_xi6_2092;
      iNsTr_162_2111 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2110_inst_req_0;
      SHL_u32_u32_2110_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2110_inst_req_1;
      SHL_u32_u32_2110_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_88",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared split operator group (89) : SHL_u32_u32_2116_inst 
    ApIntSHL_group_89: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xix_xi7_2098;
      iNsTr_163_2117 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2116_inst_req_0;
      SHL_u32_u32_2116_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2116_inst_req_1;
      SHL_u32_u32_2116_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_89",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 89
    -- shared split operator group (90) : SHL_u32_u32_2253_inst 
    ApIntSHL_group_90: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xix_xi17_2242;
      iNsTr_141_2254 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2253_inst_req_0;
      SHL_u32_u32_2253_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2253_inst_req_1;
      SHL_u32_u32_2253_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_90",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 90
    -- shared split operator group (91) : SHL_u32_u32_2349_inst 
    ApIntSHL_group_91: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xix_xi26_2326;
      iNsTr_113_2350 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2349_inst_req_0;
      SHL_u32_u32_2349_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2349_inst_req_1;
      SHL_u32_u32_2349_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_91",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : SHL_u32_u32_2442_inst 
    ApIntSHL_group_92: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi_2400;
      iNsTr_80_2443 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2442_inst_req_0;
      SHL_u32_u32_2442_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2442_inst_req_1;
      SHL_u32_u32_2442_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_92",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- shared split operator group (93) : SHL_u32_u32_2555_inst 
    ApIntSHL_group_93: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xix_xi_2537;
      iNsTr_183_2556 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2555_inst_req_0;
      SHL_u32_u32_2555_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2555_inst_req_1;
      SHL_u32_u32_2555_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_93",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared split operator group (94) : SHL_u32_u32_2561_inst 
    ApIntSHL_group_94: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xix_xi_2543;
      iNsTr_184_2562 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2561_inst_req_0;
      SHL_u32_u32_2561_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2561_inst_req_1;
      SHL_u32_u32_2561_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : SHL_u32_u32_2698_inst 
    ApIntSHL_group_95: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xix_xi_2687;
      iNsTr_157_2699 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2698_inst_req_0;
      SHL_u32_u32_2698_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2698_inst_req_1;
      SHL_u32_u32_2698_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : SHL_u32_u32_2794_inst 
    ApIntSHL_group_96: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xix_xi_2771;
      iNsTr_130_2795 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2794_inst_req_0;
      SHL_u32_u32_2794_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2794_inst_req_1;
      SHL_u32_u32_2794_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : SHL_u32_u32_2968_inst 
    ApIntSHL_group_97: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xi35_2963;
      iNsTr_118_2969 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_2968_inst_req_0;
      SHL_u32_u32_2968_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_2968_inst_req_1;
      SHL_u32_u32_2968_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : SHL_u32_u32_3038_inst 
    ApIntSHL_group_98: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= shifted_divisorx_x03x_xix_xi_3019;
      iNsTr_190_3039 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3038_inst_req_0;
      SHL_u32_u32_3038_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3038_inst_req_1;
      SHL_u32_u32_3038_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- shared split operator group (99) : SHL_u32_u32_3044_inst 
    ApIntSHL_group_99: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= curr_quotientx_x02x_xix_xi_3026;
      iNsTr_191_3045 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3044_inst_req_0;
      SHL_u32_u32_3044_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3044_inst_req_1;
      SHL_u32_u32_3044_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- shared split operator group (100) : SHL_u32_u32_3188_inst 
    ApIntSHL_group_100: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x012x_xi_3177;
      iNsTr_212_3189 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3188_inst_req_0;
      SHL_u32_u32_3188_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3188_inst_req_1;
      SHL_u32_u32_3188_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_100",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 100
    -- shared split operator group (101) : SHL_u32_u32_3273_inst 
    ApIntSHL_group_101: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= expx_x0x_xlcssax_xi_3250;
      iNsTr_206_3274 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_3273_inst_req_0;
      SHL_u32_u32_3273_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_3273_inst_req_1;
      SHL_u32_u32_3273_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : SLT_f32_u1_1737_inst 
    ApFloatUlt_group_102: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= speed_refx_x1_1711 & iNsTr_8_1730;
      iNsTr_11_1738 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_1737_inst_req_0;
      SLT_f32_u1_1737_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_1737_inst_req_1;
      SLT_f32_u1_1737_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_102",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : SLT_f32_u1_1890_inst 
    ApFloatUlt_group_103: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_33_1885;
      iNsTr_34_1891 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_1890_inst_req_0;
      SLT_f32_u1_1890_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_1890_inst_req_1;
      SLT_f32_u1_1890_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_103",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11000001101000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : SLT_f32_u1_2864_inst 
    ApFloatUlt_group_104: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_73_2859;
      iNsTr_74_2865 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_2864_inst_req_0;
      SLT_f32_u1_2864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_2864_inst_req_1;
      SLT_f32_u1_2864_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_104",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10111111100000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- shared split operator group (105) : SLT_f32_u1_2914_inst 
    ApFloatUlt_group_105: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_97_2909;
      iNsTr_98_2915 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_2914_inst_req_0;
      SLT_f32_u1_2914_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_2914_inst_req_1;
      SLT_f32_u1_2914_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_105",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 105
    -- shared split operator group (106) : SLT_f64_u1_1840_inst 
    ApFloatUlt_group_106: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_25_1835;
      iNsTr_26_1841 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_1840_inst_req_0;
      SLT_f64_u1_1840_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_1840_inst_req_1;
      SLT_f64_u1_1840_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_106",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1100000000100100000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 106
    -- shared split operator group (107) : SUB_f32_f32_2841_inst SUB_f32_f32_1814_inst 
    ApFloatSub_group_107: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 1, 1 => 1);
      -- 
    begin -- 
      data_in <= type_cast_2839_wire_constant & iNsTr_69_2836 & speed_refx_x0_1791 & iNsTr_20_1810;
      iNsTr_70_2842 <= data_out(63 downto 32);
      iNsTr_21_1815 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      reqL_unguarded(1) <= SUB_f32_f32_2841_inst_req_0;
      reqL_unguarded(0) <= SUB_f32_f32_1814_inst_req_0;
      SUB_f32_f32_2841_inst_ack_0 <= ackL_unguarded(1);
      SUB_f32_f32_1814_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= SUB_f32_f32_2841_inst_req_1;
      reqR_unguarded(0) <= SUB_f32_f32_1814_inst_req_1;
      SUB_f32_f32_2841_inst_ack_1 <= ackR_unguarded(1);
      SUB_f32_f32_1814_inst_ack_1 <= ackR_unguarded(0);
      ApFloatSub_group_107_accessRegulator_0: access_regulator_base generic map (name => "ApFloatSub_group_107_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatSub_group_107_accessRegulator_1: access_regulator_base generic map (name => "ApFloatSub_group_107_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(nreqs => 2, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatSub_group_107",
          operator_id => "ApFloatSub",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 2,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : SUB_u32_u32_2043_inst 
    ApIntSub_group_108: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_53_1980 & iNsTr_55_1992;
      iNsTr_64_2044 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2043_inst_req_0;
      SUB_u32_u32_2043_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2043_inst_req_1;
      SUB_u32_u32_2043_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : SUB_u32_u32_2163_inst 
    ApIntSub_group_109: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi3_2058 & shifted_divisorx_x0x_xlcssax_xix_xix_xi9_2141;
      iNsTr_137_2164 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2163_inst_req_0;
      SUB_u32_u32_2163_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2163_inst_req_1;
      SUB_u32_u32_2163_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : SUB_u32_u32_2322_inst 
    ApIntSub_group_110: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xix_xi23_2318 & xx_xlcssa10_2297;
      tmp26x_xix_xi24_2323 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2322_inst_req_0;
      SUB_u32_u32_2322_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2322_inst_req_1;
      SUB_u32_u32_2322_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- shared split operator group (111) : SUB_u32_u32_2488_inst 
    ApIntSub_group_111: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_77_2425 & iNsTr_79_2437;
      iNsTr_88_2489 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2488_inst_req_0;
      SUB_u32_u32_2488_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2488_inst_req_1;
      SUB_u32_u32_2488_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_111",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 111
    -- shared split operator group (112) : SUB_u32_u32_2608_inst 
    ApIntSub_group_112: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xix_xi_2503 & shifted_divisorx_x0x_xlcssax_xix_xix_xi_2586;
      iNsTr_153_2609 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2608_inst_req_0;
      SUB_u32_u32_2608_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2608_inst_req_1;
      SUB_u32_u32_2608_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_112",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 112
    -- shared split operator group (113) : SUB_u32_u32_2767_inst 
    ApIntSub_group_113: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xix_xi_2763 & xx_xlcssa5_2742;
      tmp26x_xix_xi_2768 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_2767_inst_req_0;
      SUB_u32_u32_2767_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_2767_inst_req_1;
      SUB_u32_u32_2767_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_113",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 113
    -- shared split operator group (114) : SUB_u32_u32_3092_inst 
    ApIntSub_group_114: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_x016x_xix_xi_2984 & shifted_divisorx_x0x_xlcssax_xix_xi_3069;
      iNsTr_170_3093 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3092_inst_req_0;
      SUB_u32_u32_3092_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3092_inst_req_1;
      SUB_u32_u32_3092_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_114",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 114
    -- shared split operator group (115) : SUB_u32_u32_3246_inst 
    ApIntSub_group_115: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp25x_xi_3242 & xx_xlcssa_3232;
      tmp26x_xi_3247 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_3246_inst_req_0;
      SUB_u32_u32_3246_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_3246_inst_req_1;
      SUB_u32_u32_3246_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : UGT_u32_u1_2081_inst 
    ApIntUgt_group_116: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_108_2077 & iNsTr_61_2028;
      iNsTr_109_2082 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_2081_inst_req_0;
      UGT_u32_u1_2081_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_2081_inst_req_1;
      UGT_u32_u1_2081_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : UGT_u32_u1_2526_inst 
    ApIntUgt_group_117: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_125_2522 & iNsTr_85_2473;
      iNsTr_126_2527 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_2526_inst_req_0;
      UGT_u32_u1_2526_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_2526_inst_req_1;
      UGT_u32_u1_2526_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : UGT_u32_u1_3008_inst 
    ApIntUgt_group_118: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_146_3003;
      iNsTr_147_3009 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u32_u1_3008_inst_req_0;
      UGT_u32_u1_3008_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u32_u1_3008_inst_req_1;
      UGT_u32_u1_3008_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000011001111010000011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : ULT_u32_u1_2121_inst 
    ApIntUlt_group_119: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_162_2111 & iNsTr_108_2077;
      iNsTr_164_2122 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2121_inst_req_0;
      ULT_u32_u1_2121_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2121_inst_req_1;
      ULT_u32_u1_2121_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : ULT_u32_u1_2168_inst 
    ApIntUlt_group_120: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_137_2164 & iNsTr_61_2028;
      iNsTr_138_2169 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2168_inst_req_0;
      ULT_u32_u1_2168_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2168_inst_req_1;
      ULT_u32_u1_2168_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- shared split operator group (121) : ULT_u32_u1_2566_inst 
    ApIntUlt_group_121: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_183_2556 & iNsTr_125_2522;
      iNsTr_185_2567 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2566_inst_req_0;
      ULT_u32_u1_2566_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2566_inst_req_1;
      ULT_u32_u1_2566_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_121",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 121
    -- shared split operator group (122) : ULT_u32_u1_2613_inst 
    ApIntUlt_group_122: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_153_2609 & iNsTr_85_2473;
      iNsTr_154_2614 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_2613_inst_req_0;
      ULT_u32_u1_2613_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_2613_inst_req_1;
      ULT_u32_u1_2613_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : ULT_u32_u1_3049_inst 
    ApIntUlt_group_123: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_190_3039 & iNsTr_146_3003;
      iNsTr_192_3050 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3049_inst_req_0;
      ULT_u32_u1_3049_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3049_inst_req_1;
      ULT_u32_u1_3049_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : ULT_u32_u1_3098_inst 
    ApIntUlt_group_124: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_170_3093;
      iNsTr_171_3099 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_3098_inst_req_0;
      ULT_u32_u1_3098_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_3098_inst_req_1;
      ULT_u32_u1_3098_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000011001111010000011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : XOR_u32_u32_2032_inst 
    ApIntXor_group_125: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp6x_xix_xi2_1955 & tmp10x_xix_xi1_1951;
      iNsTr_62_2033 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_2032_inst_req_0;
      XOR_u32_u32_2032_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_2032_inst_req_1;
      XOR_u32_u32_2032_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- shared split operator group (126) : XOR_u32_u32_2312_inst 
    ApIntXor_group_126: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xnotx_xi21_2307;
      tmp21x_xix_xi22_2313 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_2312_inst_req_0;
      XOR_u32_u32_2312_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_2312_inst_req_1;
      XOR_u32_u32_2312_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_126",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 126
    -- shared split operator group (127) : XOR_u32_u32_2477_inst 
    ApIntXor_group_127: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tmp10x_xix_xi_2400 & tmp6x_xix_xi2_1955;
      iNsTr_86_2478 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_2477_inst_req_0;
      XOR_u32_u32_2477_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_2477_inst_req_1;
      XOR_u32_u32_2477_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_127",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 127
    -- shared split operator group (128) : XOR_u32_u32_2757_inst 
    ApIntXor_group_128: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xnotx_xi_2752;
      tmp21x_xix_xi_2758 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_2757_inst_req_0;
      XOR_u32_u32_2757_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_2757_inst_req_1;
      XOR_u32_u32_2757_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_128",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 128
    -- shared split operator group (129) : switch_stmt_2045_select_expr_0 
    ApIntEq_group_129: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_61_2028;
      expr_2047_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2045_select_expr_0_req_0;
      switch_stmt_2045_select_expr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2045_select_expr_0_req_1;
      switch_stmt_2045_select_expr_0_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_129",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 129
    -- shared split operator group (130) : switch_stmt_2045_select_expr_1 
    ApIntEq_group_130: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_61_2028;
      expr_2050_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2045_select_expr_1_req_0;
      switch_stmt_2045_select_expr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2045_select_expr_1_req_1;
      switch_stmt_2045_select_expr_1_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_130",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 130
    -- shared split operator group (131) : switch_stmt_2490_select_expr_0 
    ApIntEq_group_131: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_85_2473;
      expr_2492_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2490_select_expr_0_req_0;
      switch_stmt_2490_select_expr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2490_select_expr_0_req_1;
      switch_stmt_2490_select_expr_0_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_131",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 131
    -- shared split operator group (132) : switch_stmt_2490_select_expr_1 
    ApIntEq_group_132: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_85_2473;
      expr_2495_wire_constant_cmp <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= switch_stmt_2490_select_expr_1_req_0;
      switch_stmt_2490_select_expr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= switch_stmt_2490_select_expr_1_req_1;
      switch_stmt_2490_select_expr_1_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_132",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 132
    -- shared split operator group (133) : type_cast_1749_inst 
    ApFloatResize_group_133: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= speed_refx_x1_1711;
      iNsTr_13_1750 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_1749_inst_req_0;
      type_cast_1749_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_1749_inst_req_1;
      type_cast_1749_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_133",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 133
    -- shared split operator group (134) : type_cast_1759_inst 
    ApFloatResize_group_134: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_14_1756;
      iNsTr_15_1760 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_1759_inst_req_0;
      type_cast_1759_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_1759_inst_req_1;
      type_cast_1759_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_134",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 8, 
          output_mantissa_width => 23, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 134
    -- shared split operator group (135) : type_cast_1777_inst 
    ApFloatResize_group_135: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= speed_refx_x1_1711;
      iNsTr_28_1778 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_1777_inst_req_0;
      type_cast_1777_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_1777_inst_req_1;
      type_cast_1777_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_135",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 135
    -- shared split operator group (136) : type_cast_1787_inst 
    ApFloatResize_group_136: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_29_1784;
      iNsTr_30_1788 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_1787_inst_req_0;
      type_cast_1787_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_1787_inst_req_1;
      type_cast_1787_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_136",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 8, 
          output_mantissa_width => 23, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 136
    -- shared split operator group (137) : type_cast_1834_inst 
    ApFloatResize_group_137: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_24_1831;
      iNsTr_25_1835 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_1834_inst_req_0;
      type_cast_1834_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_1834_inst_req_1;
      type_cast_1834_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatResize",
          name => "ApFloatResize_group_137",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 137
    -- shared split operator group (138) : type_cast_2215_inst 
    ApIntToApIntSigned_group_138: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi14_2194;
      type_cast_2215_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2215_inst_req_0;
      type_cast_2215_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2215_inst_req_1;
      type_cast_2215_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_138",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 138
    -- shared split operator group (139) : type_cast_2269_inst 
    ApIntToApIntSigned_group_139: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_141_2254;
      type_cast_2269_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2269_inst_req_0;
      type_cast_2269_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2269_inst_req_1;
      type_cast_2269_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_139",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 139
    -- shared split operator group (140) : type_cast_2660_inst 
    ApIntToApIntSigned_group_140: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= tempx_x0x_xphx_xix_xi_2639;
      type_cast_2660_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2660_inst_req_0;
      type_cast_2660_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2660_inst_req_1;
      type_cast_2660_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_140",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 140
    -- shared split operator group (141) : type_cast_2714_inst 
    ApIntToApIntSigned_group_141: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_157_2699;
      type_cast_2714_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2714_inst_req_0;
      type_cast_2714_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2714_inst_req_1;
      type_cast_2714_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_141",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 141
    -- shared split operator group (142) : type_cast_3150_inst 
    ApIntToApIntSigned_group_142: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= xx_xlcssa4_3107;
      type_cast_3150_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3150_inst_req_0;
      type_cast_3150_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3150_inst_req_1;
      type_cast_3150_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_142",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 142
    -- shared split operator group (143) : type_cast_3204_inst 
    ApIntToApIntSigned_group_143: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 1);
      -- 
    begin -- 
      data_in <= iNsTr_212_3189;
      type_cast_3204_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_3204_inst_req_0;
      type_cast_3204_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_3204_inst_req_1;
      type_cast_3204_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unguarded;
      reqR <= reqR_unguarded;
      ackL_unguarded <= ackL;
      ackR_unguarded <= ackR;
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_143",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 143
    -- shared inport operator group (0) : RPIPE_in_data_1720_inst RPIPE_in_data_1723_inst RPIPE_in_data_1726_inst RPIPE_in_data_1729_inst RPIPE_in_data_1732_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(159 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 4 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1, 4 => 1);
      -- 
    begin -- 
      reqL_unguarded(4) <= RPIPE_in_data_1720_inst_req_0;
      reqL_unguarded(3) <= RPIPE_in_data_1723_inst_req_0;
      reqL_unguarded(2) <= RPIPE_in_data_1726_inst_req_0;
      reqL_unguarded(1) <= RPIPE_in_data_1729_inst_req_0;
      reqL_unguarded(0) <= RPIPE_in_data_1732_inst_req_0;
      RPIPE_in_data_1720_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_in_data_1723_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_in_data_1726_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_in_data_1729_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_in_data_1732_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= RPIPE_in_data_1720_inst_req_1;
      reqR_unguarded(3) <= RPIPE_in_data_1723_inst_req_1;
      reqR_unguarded(2) <= RPIPE_in_data_1726_inst_req_1;
      reqR_unguarded(1) <= RPIPE_in_data_1729_inst_req_1;
      reqR_unguarded(0) <= RPIPE_in_data_1732_inst_req_1;
      RPIPE_in_data_1720_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_in_data_1723_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_in_data_1726_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_in_data_1729_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_in_data_1732_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 5, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      iNsTr_2_1721 <= data_out(159 downto 128);
      iNsTr_4_1724 <= data_out(127 downto 96);
      iNsTr_6_1727 <= data_out(95 downto 64);
      iNsTr_8_1730 <= data_out(63 downto 32);
      iNsTr_10_1733 <= data_out(31 downto 0);
      in_data_read_0: InputPortFullRate -- 
        generic map ( name => "in_data_read_0", data_width => 32,  num_reqs => 5,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_out_data_3305_inst WPIPE_out_data_3308_inst WPIPE_out_data_3311_inst WPIPE_out_data_3314_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 1, 1 => 1, 2 => 1, 3 => 1);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_out_data_3305_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_out_data_3308_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_out_data_3311_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_out_data_3314_inst_req_0;
      WPIPE_out_data_3305_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_out_data_3308_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_out_data_3311_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_out_data_3314_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_out_data_3305_inst_req_1;
      update_req_unguarded(2) <= WPIPE_out_data_3308_inst_req_1;
      update_req_unguarded(1) <= WPIPE_out_data_3311_inst_req_1;
      update_req_unguarded(0) <= WPIPE_out_data_3314_inst_req_1;
      WPIPE_out_data_3305_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_out_data_3308_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_out_data_3311_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_out_data_3314_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 4, buffering => guardBuffering, use_guards => guardFlags) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_173_3297 & iNsTr_67_2818 & iNsTr_49_2396 & iNsTr_39_1941;
      out_data_write_0: OutputPortFullRate -- 
        generic map ( name => "out_data", data_width => 32, num_reqs => 4, input_buffering => inBUFs, no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- declarations related to module vector_control_daemon
  component vector_control_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module vector_control_daemon
  signal vector_control_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal vector_control_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal vector_control_daemon_start_req : std_logic;
  signal vector_control_daemon_start_ack : std_logic;
  signal vector_control_daemon_fin_req   : std_logic;
  signal vector_control_daemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module vector_control_daemon
  vector_control_daemon_instance:vector_control_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => vector_control_daemon_start_req,
      start_ack => vector_control_daemon_start_ack,
      fin_req => vector_control_daemon_fin_req,
      fin_ack => vector_control_daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(31 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(31 downto 0),
      tag_in => vector_control_daemon_tag_in,
      tag_out => vector_control_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  vector_control_daemon_tag_in <= (others => '0');
  vector_control_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => vector_control_daemon_start_req, start_ack => vector_control_daemon_start_ack,  fin_req => vector_control_daemon_fin_req,  fin_ack => vector_control_daemon_fin_ack);
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end Default;
